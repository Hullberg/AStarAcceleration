��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���q�����W�E�9 Vοօ�̷�S�;(B�����",�U�s����6���i	t̂9։l��cE���	����a����	YD����>v��<�b����)a�������⚴�i��A�Z��1�С2�1��V��@��zM��՟"Zq�~���aˋ��I᭗6�����n�k�a=,�؆�A��O��X)j��Y�>]Mu�v��B�.F:R�c���5��v������KU�;�U���H�
�l��'�K4�}4�c"jcx�nOd�F{��Mf�['>[���B�a�r�>;�~���1��8�W�8��_̀Ǌpz!n�ʑ��<�5�Z{Y�?���:R��-�{8{H�
�pM_]" R���%�I�8����ڱJ�!vzoE��}GP�����4_K��t�_���K�����B������g�Y�����������b�<���65:s���c��X�[��QG�77��^!�x�*��bU�=ȑ1��(:��^:R[�@�,���3�MTC���"�h(EJ�;lς�]%����J���
���+|��I9��W$���UT��yޯ#�E.e2��)�vŅ�]�1���1���:�'Ua?� �x��i^�u٘�m�+Ŏ��j��S��B��<�/\͈�6���Ѽ�8�b�uQu����(#(m�/�XY�X1����Ƅ����1~��F	sq㐶*m�� �G��Mj�=�Qhn��d�+R��m��˥�vZ�����8���1�E���n�/9��f&C��G罵j"ү�fϴ��<բ���x
O�:u_��v�ze�WNӥ�W6�y��J$�	2�/�v[c>��e��yoŏ G6>'ŝ_J���YN�hk�W䘐��8MmqSФ�pk������U0��vM�j'�R�5c�,���1`���XS����	�!�Î�@/�)W\�Z�nB�B܆�����ϔ�H e��Q����5��v^��)ź�Fx�'ߞ�Em~A\���� m�?�,�F/��7��!|��4goN}Ee���/+i�ouMY��&+톮���~{�'�����2_ʿ�t+Vym� @����u[�C3����2�c�|���{7�2(�c�l�73�˭�ώ�9=��g��A㊪��d�#���F*�ѥz���E��鑦��%��8�����6	����]�D9�C��}tsb|�#�,��\�M�c����xcڅ(��D@Ȱ[��WR�lTѰ��H��F�٨���c���Y2�z�1yIՉB�e�0�,��no2�0Z�2)D=�?�_^������(�)�H�H�*[My�W�)��S�Z�z�k��,��<�'��v�.��|��R��8�����\�Y�/M�~L�zc#"��F0��%v%�����'<_K�rk��e�����Q̳6y���6܍�W,	Q����K\�4��g��y⃯c>1$Y�~�Z�wt�'%�noh���t8Q;�J��1ɣ�+6�F%s�����i	�l-�Zs�iio���T�G\�0=��-<��@rJ�� ȏ������ ��I�r紺��eJ���flk~���~|�A=1ᵁ�}�	-��'���=#�� �-�>�[�pX���G��$��4�QJD�bA�9�b%b�"��1�A�-ϙ5y�sm�Y��I+��.ksu���^�t��^��{���w+�`�?����*����N�/���W�șG�:�4$| h!���3�ˌ�^�M'z��v\�F�v~� @rSUΓ�DL�wk���<$�^M֍.�v��{� �*45�8d��Z�_I|��e֐��Wvt�{�˭t%��8���c�:5��Tn�1���pD�T�9��٠J$��i�^i�,���,���B2#��=�4����}��N���-���U�5��2�RBuS��K�{�Ej͂��Q=W���{k�R��Tr��p�-�I�/�.Z���:�zeo���_�F:�F��N���U��}�<��`0@��vYT�J��7*{�<�}~Ҡa�.�:E8�I�9q�y���E� ��!)�)vT��ǡ�r	����0���C�-W�kw�z+J�ۑb�5G��9�zA��S����0��!�o[R6�Z��Ѓ��U/f�e+h�Ş=���b0Sv�
�g���$;�|���kV}��F�ò�S:o��$d5��>��V.�5��Q��\Hm��"'tj�x�8�E��X�~�-6�;棕�3�-�g�_1/ff��i�Jj�ux@����t������O�7wuM��=r��	6�������8�ߐ��|cW�r��sD�DVN�ʝ)/��^["
���u��oRH-�Ҵ��D
��C�+���c��%��<QC�����R[ڝV�@������1%�x���5ˬ�ߍ��R��w3�t�ê��%��>UQSJ���H�Q��{w$c�៦�?ؖ7?q�f��ix?��[!���3nws��]�GP1&���In� �[��9�lq�g�\N��j�"̆RO���O�#�r�%�Vhغ�TN�K
�f"�ȬN�)`���R8�����&�������i��'�`P�:��9�Վ�n8�x��nk�m,�����V��/ߖ�?�O[�2"ʷ�Vß�˖:+_���{	�4�G�޾F߳9�z�(U5T���07m�����@<$�������o�{�e��EB�;�*2y����D�Uշ��$�'�.v15"����O�qK	d��$pc¿���R�+9Z��E�
X�2�{����e[�r|��4�aB	Rg��=����g���1迉h�*5q������(�{��ȇ�\��M��u�e=�kt�D@	-/;��S4�k_\�[7���z�B����F#�����g{��9���Vj#^�Y�9��������q#��ox{w�b��fe��^����� �/a�"ƣwnB���{h�{y��B��Xi����~�����Ǣ|�U�M_�G��0㝫�Y�`�S�?������9-�}x'���.���`.����6�"O��O��:� gw��N��)�4tlԃ��޹�1��u�����H�,�Ó2n�?��-BN�-��>��=��pd�𱰖"׃�2�9޶�F%{��Ғ���ٓ��#��yXF��F���E���?����r�PP^,���H��8(kV<���;j�jm)�R��s��N���*I�%)?ɖ��˧��-�d��������#��I�N+Ȳ����8!g�ڠ��*�C̄�;���ؒ�1�xl�(�����.�� lt%E�HNE-��g�2k4�s�[O���IPX�.��ҴK��:~�S�����6D���gY&�4f������۳Yo을��)B������=��$����
�yPt9��yZU���n/��^GZ�
q��+��O34)*������d��U�ʛ�:�9ZX/p45���~���T��1
^�#���3
�A������0q����ъ+�)1��=/b5%�?H�ͩ �z�(��2����DN,�G?光�����2���m���wdGw��ҧS5�|�]o�8&i^pI_�R���@�d�_�s�}�/L�(M�JP�k���k�^\q�Y���4�yl�	��o�DTYe�j���^]�ϳ� �ߩ"�1�L-u�k�S�1E:ݞ��5S{�����9��B�{Ƃ�ڗ�گLj)8�+~8���?Rm��SYH.񻱕/"�bO�o�m���T3D���x�9�u�r :�1�Qop���6OL�_`�
���a(x~�bb $cS�hzh�� ��h���y��z��G-z_<�=Wa��è�Ԭ^��X���V%J����S ��%�����ɵ�
�WFs�_�j��AE���9��\��b�o��-C]щ���;��~?=ԏ�>wh	q��L�AJ ����%i���	�ϔ��Dn�zBC �5s^�:��",���[��ʋ]2�'�ܗ���
��<YHva�V��,��^� t�������N�� �S��H�Z�g�wS��Wc�w���S�R8΀{S@���Ƞ�M�Si��;�k
��U@����k�
�<]�w*��B���.
��IQ9l�aX��3�+nBD�Z� zM�`�d�=t���f<��B-	����7��8x�P
�S�)
;)���Ѽ��"���=���,+cm,y�@�������Lj��j�NF��8�Tꯐ ��OV��Q]��z+>KĵtW�.D~]���-��t[!�F�;���j�;��v�ݩ������S;IVêC�
�]qO����iY/���uT�4�H3��AjGQD�9}p�R/n�&�l�C��	A�spW�!�̳)�K�����c�f�-�b1qT�ϱ?�0��)
ZX��������/t
�/F���4��B����$�B��P
��ޒu�A�Jm��=����\�+H�* �c��L7>,4���>����t��4�E�_�8F��7q��<=��!�FyKë$>�Z�]�	'+ɸ�/劇�S��%�W���������4�}+�����ޫkX�T��N�f]F��Bv�9N�3{�2�Y���˻����3�w\�py������ˆ�~���^Z����w�`u���@�E#?�#2��A@p�"l����"�I���~�R톜�Z�'5~ nǳh��+
��>{�dy��L�2�5ޠ@�\S���h�j����χt�
�c njث��B��b�����	�1/�T������	���$�K�aKB	��2M����8ھ��7�jIA�kp!����a+�F�Kٿ1>���Iz J���1�R���J���"�!���*�dV�2¢y��_8��Y��z� H�>_�r��j�%�����풆���XG�5"W�c^�JԲ���������q��.��:K��N�d+~�?ț���:�·�
�)6u��D�0�~�zv.>0��pu/,Ͷ,��_}ԍ���CQD�'����Sc�P'�m��D��y�ͅ�Ff8���yo����1Ź(e�#����4�M�"gXn��H��ȥ@֤�]'8���5*�g����/�S�?9(�K���BǶ{�w�G�q@�7�ο�8�
�4Hm�%���a�k��	[Ŝetr5^�>W���p������cbχNjϱı3�H������0�XA��oe��T�{;��e�2&jY���5H�1㏜���9��UWAQ�3� �0��0���"���&�b}������+�Iǋe睫	��a��yD�3䐨�'��$VnZ�K@����0���F�U���;[kx���)�cG���/d�]�d�&�eWi�g�{�x}	�|c�8��Q~�(mM�q,sQ���x��uxf���5^ 9��
��m�w��z��z9rT�=�W���$ƪ�.Ϡ`ř�>1l@L쇊� �C^p|ߢ�����ֈ�&��fq��l�痚�?���i`Vd<aNh��H�,��6A{x�b���1o�$�w[C�5m�:�������!E�\U�L^LK�
I�y_�u�m�<�N���0�8�K]�������V��eG���<��>�2��V�#��^�h�k&�ڢ쪃�7��"Z�p|n�@���� ~XRڲ�զ�
Ҷd�!s�������	�{�:&��C,z }�z���4��al_E����r0�d���Rg��t�ձ:�Ƭ�9��e��q���ߊ�t�3�|�[���"����,�R���}s"���@��p�xJ������S�xf)���F"��1�W��͟u��23��P�f�vn�B�u�{� �|'C�`rN
�WV���3��Y ��5�^���d��%�=�[Y)`���k�jg���פ@f�#6�K�;d�S1s�M��k	��6�C�3�B]�.��d����!�D�� ����K�-/��zd��񞊫*4s�]V屑<2�EQɘ!�V�:�8��%�UJ� �e����NT��'f"3?�\�P :k@�f��4"<D��,�ʀ���c�F);1��Zuu��$�-Un`�>{fܸ�X�8���2�Z��|�Ƃ�C�����4�U�&�6>��:�0	��f
m�nbs n��RR�s���!D��=gc��Ԇ���N���1pQ�����A�zw!�N�_4�rڶ�N�c�_��ܚ�?�y��-}��\헐�s��k��27LV�5����򅬩�5)���i�ְ^��ْ����.L°|�EX�4���������bh��t�G�|H�Vj��Ek�Zx��<c�S��B�b#ܧ<Dӯ����'��*1q6|��d����a�>31}{L]�	Ey+d����!ݒ:���u?7e��l$WBw�9��U
�-j8"�e]�RR3��T��]� C��t���F���*��|W��/��})���K�Hn�=���0�x��Y�6K��l�P�pda^[��J%Nj?{�B��j�92�Kt���5piEcP�E�>��YS��X�V���b�J1���?�{�
�uPd`��X������4�E�d�{����iHe�;��s-V��:�X�0eJ=��Iw�� E�.`�� U�9�M��|8˵����b��A>2�|模ذߐ��d,s!fӰum�l��sP�gs����t�
���c�f���˫�SԜ#���k������#�'`wi��T�8�,H4�@���ܬ\���_<�s��-�{�7����Z�s�3��$���l6�9�AQ���� *8=%OQ6t֩`��;	��,Vx�tb[�b���>�K��B�$U.U��#�4�����g��y]tI&�x'�5h-x��3��֖�LI������sxJ�U~{����\�a����N^f���i\��2����	�}����RhBf�Sޱ����]����\�V����+W��Rϯ��E���y�f�3
Q�Gf�Xp�ԥ��Tg�_>�ǯ�@(}� +��^-�S4���E=O�R_+�<��`1�1��֔��b��xP����'̂�����������8ӭ�A+����;�:w8{��>�l�?(��q��Hܝ!j�X��`�R�E="�'Y�HAa+,NC���W�y�ǐZ��f�u� ���F�6n��Z�{2v'G���wj��PBz!�qE�{zҦ9B�=bp{L�[�������=Jpn�k���%ֵ���|�+'$A	j�ѹʵ�2�ړQ�LM�x��3��2Kr�&�]�/0� �)?b#.��������|����]�ՙ�-*ю[��c�V��oK*$�Pff�\�u�C�y89��<~�끱���$���j� ��o�U�#��Bx׻^'gNԳ����ꙀX�K���L�n�}��{{6m�G̟� dQ=8�P�1�{�R��_�V� �(�Z�<!����da(��2�����nzI�'ǭ���F7C�g���� �����}xs����`=G���6���H�r�Y ��������R�baL�$RȬ�����P-@���<��A��(.��c@�z����<7��{���Z�2)�/���[Ʉ\�$U<�Ĝ�<^�b��ӯ.�O_�;%���7��˨]��%�|�8Q�����f�����$=�uoW9(ǳ$�q�����D�5��R��(P��:%��A!>�����1"�c�v���t;v� n�`�yrd�t���֟|��K=���n���鵟�b�G>Ȭ#7}9�����O�St\?���m��&v����mC��OT>b�iW�6� Qj64��Qw�p�G����:�hȈS�6�Ը���Q0�#��vKy�MO�x$�8�-#���Ɇ���l=��7M��R�%a�N�ŤpW�[���`i`k�x�)Q;F��qhD1�y�<���"Nڬ7#��wAD���e,�E�mm)��l�u`u�%ۃu�������du���N�	.J�9�x��2&��q�cUE$�[�*P�©[��`��ɉ�[x�B�hh�7w���kl�mގ�
_~��lz���c�r6�ᓙ���D�4���vGo�nӂC�Nç�AS˸�+���ڱ���(ir�ƹ�_W����s2%�n�����eco3�g��@�l�4�t���"]�C�q)�I^�C���s�1-d���^2/d�ǽ˷�5�E��sY�� {Q��]f�q����ex7�A>	Y�M����j��=V�dBE����f]�,�,��_�Hbh��MⲌP�û��YݟA�\�w75 ��M�݋z# e�b�� ���xY�[���h��ގ89�m��&�N��a�I+k�hm��� D��T��Z��0�@scs�����X�y��y�y��ґ.�>1�jYr�V����^rSX����Z�g`���m���)�c�?U�����E�=A�"��5��Z�
.���V��L3�F�K��!�A�>*X��;ljk���F�k�h�X�?�����jjb��P~E��mD��Ȟ/<0Hz"O-U�CUAu�]U�����@Þ.W��A�J=+S�/�!	��?F��Ă8ᵯ5Ƃ���
Zs��T,V~%��Xj�u�-�ڧ���=W$@�l�h��:Y�L��+1�
��k;��o�(T�1̛�ۋaЕ!�IIS8��a�<bfG}�t��\!Ț8n�@�>��@�I*��ħ�����;l����`Z��:��o��)U�EJ��b+t+�i�T��{�F:5�7`W��֦�c�VM����:va��B޿�9 ���_�6I�f8dO�;>�����)6��G
��j�ħ�!E'yf�! `fŁ�6/�$(�m���X��������.����!]���L��SaoI#Za
ȧ�)�O�쑆mv be��ᔥh�&�w%�?�^@\V�o��_4a��@)�+)*yH$!�k�M5E���h$�x��~�-�ar�Y~�syFT��?��n����5���#ȣ_� �ڪ���n�F�uj+�P?��xlSc{�PlVw��!F��2×���
Ϫ��Zd�U(��Śѣ�aCu j��#�Hx���`pz��J�(��a��5˥�7n|l�F�$��a�A?r!��/�3�VY���! �{�X	�Ir��R2����7L3^1!N�Ƶ��TZF
�-&5��J�n�jU�Qc�.��������
�V��/>�$��&�L�wA�%Idfu�2��=��b��D�^F��[2���`��5�76L�,�j�R�s�bd���n=��H��N�9���~^pYSM�=n�e¼Y�F�NX�$�� *������<�e�.��-���Ͻ��6#L~�8k����Y�|Dq�u��V�9��@1����K�/mW��y �@�T�<Y��N�cfs�C��i#���6�0���Q*y̚y+�I�Oՙ_1z�(7��*g��NP�e]�+V-"����i�T�G��7P=�&2�j;Z�e}��0"�ز2���L���ƍ`t��ܲ�v\9�_��#[̦�O�Ij�"PŅ���ď�|^��Ӥ%�[�5��>*��Ws���"d��-rX���I)b�E��.���0�J���}�n���Q�����Qҳ��|��8���M2�T�[�>����J����pD'm>����y�x!��"�`������xY� ��x�`��󂖫&\D}Kh1�[�j.	�$,�Cbp�O��=�t�����YxǾ�������@��#�{�X ��{ze�k[=�
�ɨ�A,�	
0C��
��g>(��Ӊ)y�UES�K&��p�>�9!�k��s�^���V�S\]Ƽ"Sإ��-�b�ΐ��A\��j���d����WR{a�ꡕ�i���;��0y���:ea��o��o�y	�FA"�c\����1o�p��G�SH1۾Ũ���tx5������
�|��Sn�*ߚ��Ћ����[�/()���� �u��O�b���"��~��/�t�0��+�����=Α���=^�(LC�*���W��̃w��|9�,������3��kU��s,��q'1�J��@��/e~B��&iq��%�B�b�e�����q�Dr�R%��1�g�3p����-mh����}�S�n�b8n��iGtۜ��?�|,E�_�����9T-��9M��Y��e��s�]�en�Ϝ�%���\�7�0�X�n*؛c�;ҙeXX�� ����NB�ρO��	[că��H=�0�����A�,�f���"N	�=7c|��k�
;d����W)��}3����ܐ��d�:u��<A#�.�N�Ou���Sr�����w�l ��]��� �αW�烳�'b�Q\15=oS�f%�'�"{kBnɲg$T�?-k�ېEm���[���
_ꁘ� қ�����Y(�WQ�d,2fx:Y��d��
N�^qE�^gZ�EX@p�i����hE�S,f�v�-L�V��f�`����2=GKJ�#�\�+y %1X���y���=�Q�}��|� X�GK:�����؉��u��5�'���Dvj��������Z^�!�~�&�D�����q�R��:��F�s�X�����Fa�a�6�g����p�d&��T��x0�uzHj��J.�0���;�X�V����Q�Fy{����p|i��&��Li�^O+�j3�㷐͋��3�%���:�Q�
�����Ts^wڏ�#x�����(�w��tCK6�����R-o��2�_3�E�_@!ս�K�J��+i��ŐT����T��i⇧��zd�QHaN`e�d"37���-�h�g�ZHH&X/�m�B]�^`�$�!v����!�C���4Bn�r��r�Q�:��x�_[X*>J�{�}U��[�4�l��ul0