��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���q�����W�E�9 Vοօ�̷�S�;(B�����",�U�s����6���i	t̂9։lo���M�"2s���i��훳YO����g����_�V[�}��hBNՏ��W�����V�l0iNS��?��tN�:��/��Q�y���C?`�diB�݂�'��S�BM�������
J��FiR0qvG�)穔�F}��y�`�_.^o��0A�v>��(��le�j�Ӛ���UҼ� ��!�$���tM=�NH}&����ec��ōO����K줫��,�5sAn�'M	ʈ�8*�NS�e�x��{�����IP��ԑ/�4���B��`jxZ��(�ն�d�_UK�8�����P󿨑�'$*��^Y�KT"{C�H�Uqoaѳz,譆lT�HjD���뺇����]M�e)�9�գ�$]��Fp?�&��������.���|F��u���5������P�?p�:Oym������	���T��?=�v�灱ȷ���I�4��m�'*���FeM��(?���S�R������n����*d�� �Y�18ļaj+��8�T���W�N�BT�Zӗ�8���Bz���&�숗a�������~(��H�?�&w�.na�.�ڛ��GP�s��'Q��}�Ȫ~���$�n�ü�����P:��.�3u���Ay	#�ǢZGjg�,�t�^-��R���%^è��S�� �A߶7��x83������;��6��)�B �i~ș��$�H�7��^lI<	%��)ж��$u���ËJ΂U�`���Q�?X+5���
��jl:������!��n�!�ϟ+��.��E��ʽ&�h�����D����dU���l݃�%c�%��8�to!� D/���NZG�A6�Ip{�3v���Bc�rf1�:�P@ls�$X�,"t��є�(ok�t�<�y�����U�^�nl#w���,��p��A�O||�	�%��;�٤��H�xS*꠫vb��5ٛ=���#'��/(���cWZ_Y�:}(B;	5M�@��޹�/�-�p-ǟT��#��`���y&��d�<D�!���G)0M�5�U ^���IyL�h��o���< ��<=�aE�]�:u��vB� �졥�c�,���A(��P�C��l�W�*Ct�\"%l�J�)A7�K�Ђ�1F������������h�^pIT�X��8�ڿN]��|}2\��;�~��HO��$�Qu��^�B2�[�0Q�ؒun����¡lVC��j��ҹ ��y\u��{��#����CV�{5&TO�{�F���k�ewi�ԝq��Jh�8���-@1=�e �y�lr�ٝ��� �f�4��d�|�wɒ-���(������uY���U*5F�Tnp�P���}���b��1�
�4�X,�<#�̙��4{	!��#W5o�]���Υ��f���fjƲ$��K8�-*��As2���H��P ^HA62�@!�6��z�א� "c�	-k{��t���Q���p�E��4��X�Y���ö>+��j!c7�붗}����ͭ�#�^ �纷�q�R����]�BDh��}O�g������![^@04Q����F�"�s��ZɎ��e��(`>V.U���@�JӇ�b��ݙ:JD	rmt�Gj��B}�)�Jl���x�^<8�7���}� ��jK,0����s�yʙ{tH6��[r7�ixΐ�e�ëߚ��T��V��xۂ��]�`MQߢ-��7$�TyYs���f/lnB�)��������P�y��5�-1-� ��uM���Gy;v�z�U�?D�
��D��=zq�I��a]��7���cd�TC�*h�M�+%���$O��;?%���$��"QB��������C/ts>P	dSX�s���,� %���җ��޼�#^fT2ܔv���@\��ê]V����� �Y��h����?|���n��|���Q�R���75L�
��Kأ0?}qf�L�W�K��@�1�{��Ɵ%�r�^<?���w�^�W/h����B���G��ż$*��O5�(t �-�\��n�OԗI��f�40�����C�f���۶,>��Pf@��-)ϙ��知R0�"x�6���;�������(Ls�E(���eB|�Ȃ1[�ί,p���^����׹��ZT)��j�O�G�w��v�� �X��c�j��=슞6h�������nￃ���5�(M�&�aHr�k��n��䔽g���5������I��V|<mǚ�Nl���T���8�a�7��"��3;�⁒����3��'����<'�_�~"���� .1�R��I=1�
�m�)�v�g�Ke�2E{����M��w����Tx�"0H�6�'&��F8�������/x�ߋ4�X�9��yN({�5��vB�
��e1q�&

�ү4���Vx�(R����R2ܖ3e%�^�q����� �P��{A����o¶�����G������L<;y�K�4ktm�ÓnW56�����ɤ�O>����E���ӊ}� +��	Q�Ħa^�W>��6#n�xS)	v�'Ff���&,4�Mf�5���i+e(�ٱxt�=�^o9�+�������҂�3H���+-Se��S�+��x�������9����v�ě��a7_]i����M����05j5wVQ2������g�OX6MQ���>�:_��2��哾7aʑS�Ri�60$kK����=U�Ix�u����>&���79$@�Z��mL��0J���ы\�&�,�p�:�k�vt�Yc��wr^��&א������/֭F�󾥛`���\v$��/��_�$ 얐2�����z��>%�� &��ֺF�[�G��Cq)DP8.��L5)K���j�|��I���о�u�Y�&/DF��b�x�0��Q�;߶l,�M8T�Kqqs�S�s~fG7_yhwu\S\�o{��E��q�����}���F��H���L��h��"+�&Z��{�}����w�����1"�${�;)a�� �7�C����-���x0�nGw>�7Y���^-qs�gA��q8\Ex`eLE�x~/y,W������q])@|I�S� ��g4��mp6M����\��6wy�:�6���v,���7q�+!I�#�����A*g.KT��(��]0^z��+�Z��4���+��{�C��UlIE�pS�������RE�pv�a�A�$1�5�g��82w��fs7z�����f��h�78o�cx�/1+��~rdU�~C�ͩtVI�����-�(�w}�G��I���$tf
�Mn��V�0�yi;��rȪ� >�ρ�~o?��G�&��jMpOT�LJC��#
Hu�q�d���'��L���5YzD༬�<���	4��ڇ1���Qe\n3ơ�\���_��ً���w�&R[��pQ� �I��o	T�}ȋ�Uȍ���D݃8F���||�Z�Vr/� �0�%L�,~ę��zg�)����<��x�}�U�	U����O�I������Q��zu5V����!׽�U�]��
h�-�
'*�'���7���6_��竕E2&I�f��]�_�j*2ץp��Z�9F���T���4��������-�(�n�!6��m/���!�Cq,lY��RL��8����'0%��U:ry?���_n/榇���
�%�"��4�TT��Oʷ�z��>�I��b�&]�t�~�~�������!�Y�)�\�
�y#�D�w����J>ɛr��#��O�c|	��]6AX�����0�
�_Z�]~z��'��!��U��Q���lr�ᪿX�طV �⦑@fsc���B���g��H�g}f����%�{CY��:^y����`�A�d�8�����C�F��#q�������/�)O�y���j8�2k��V��^��縃��iYަ�q�c�H���Cψ9�(�?.�V�1^+σ�Mн�t�7'��t�
�8�mJٻ40��#���'��
�l�d��j�ɿ�ǙS���	C�P����hUz����5�WW�&i#.)�`CG,`���$H��|�UI06��sI��_��v)K	a��LV�nȶ|���6�G���������y�������Zh�_EsJ����쇊�0~�XK�%8�\,p$��wl�/�
�L��m��xP��d���o�8��m���	?�{|��\��*I��=s/:f 8��nF��U��RN!�ՍsI|fA+���=�T���rl=��s����=ȭ�_ �W��kׄƟh����ƕ>5yn�L�����hj�@̦C�Cy |2,��`�����.��Eo�/����0\2RD
TFaYF+����5�=w����9$�Q�;;���,Cʚ��t2�B�|8xA[���h����t^�T�z9�/�F>��
�tgOqo�Aw�����fW=D`s��(���N�}�i���HjgYj&D�����+���?�V�k���4�_���cؘ块?���h	7��[�Y	�7t��$���[�`�u39�PZ�?���4���6�:���8s۾�z�2o�_]� ���
�6�y�L��t��!�|y�o���w@3䟳!��@�P���+t�<"Z��9�1q�*���(L1��j*_�d�\Ot�ʰ�J�吷x�S�*0א�PI���\wCa�#�y�n���(���r�6S��]���D�d�m� ��'� O�ΰ�I :��t���<���#Ƅ�K
.;�y�[q�1�j!E�������cư6�kB�݆ܚd81���G��t�]u4�^p�qr�Ir��o�uVD}kJ�̰���sq#	-9M@�@[�2�j��IQ��ZA��Jo�H�V����**bn��߸�k�c���^�/�R`�S�iM�+ ���Z ]X��d�'[1���[��$��F׏�1Qݸ��?L�(c3���h�Q��m0�I�]Cʔp�~���>������)�^u�}�	K�	�7)�c�����~��Xi;��ۛu��J�2ܵ�dT���5���#���2�3j�0V�Y�t��!�(!rN�}^P��S۴0bٲh��Y�������D�p6i{�~+a�rLw����d�5��K�e��M:L�nT�r!�;rsR��M������:��0�\�!����4ڑn�:�Qj�ό%w��5�()ķ�dL�����P�:
�'۽v.rV��"��s~Y-#��7�ʭ.

ۃ�~��{B��9^I֒G��ϏG�W�I�;�׏Ԓ�049�t��0m�^�I����5đ�M�:�O�!�p���S���ۇ�)꒫|�H$�'��}!�$E�M�X}�J���<Bj۩� }�SaVňI��}ImmF������1�i'?��B�	@�5G�Wz2T����<���
�*Rt�b&�V;F�5�����=m�/��y���Á0a@C�q�2VR�_�T������e�P��Y��T�s�qN�$4hbs�.o��v�E���):�̶:�8�xcª70Z���_+4%,��ضn`fT��.���=��ҟ_�b[�#mh���OK�][Ȃި�Hp'( �!��ܷ���Ei�L��$oM��G"4 ��*��&��RJ;�`�V�8��quk���-�:��~=���d��L-I1=}JaH2�0����Y�$�d�����?!��K(�gJ�{���ꭾ'�^�2?���F�/������B�c[�R�|h�s�v��b�t�����;���7e���?�w��σR�!H�E��}u��`V�t}k�%��=E�Ѿ1$w}X^�K��U���)!������Zb�� ��Lߞ�,�}@��=�Fw��_�#h
�W���b|o^%�pi=����$xN��)����?<m�w5�P̬���h�!p)�Ȼ�6��MA�� �dǕe螝��O}H��3$.l@���ɑ��1��y��F<>���Qq"@ܹ�9b����~o�U��g��4.�䋝��yD�E*>���.݈s���#����#~�_]���w���3��2I�)�����%-2�&8Q��*i�A��b7�����R�r�e+�AD��2�U�U����4V/�c9s��P�ӆ�)��v� ����t�E�~�q�aS��Y��E<�.���4oٺ�R^��yZ�Û�9Ci&����þ��,b"ZS8�$Z�.^�E�4~��r���Īn��bg!���H�_��� �4��@P�5���v$��76�F�'r�M��+׎�����ɇt:�<��0"a�cvdp����w��*`g,ӥ��1����sM�Af^Y96^I(� �;3�t\]�$6���e�����\8] $H@kώ�����SEX��!!ye�����e���P!�%٥��oT�h[>��
��k�A��,O�Wt��:�u�:��-���H3�I{Fo�=����q�����P{�3���ʔ�ImY�n�t�=����o~�h!G+����HwA��^{p!ŖF&�3�1�X����s��z��9$JG��� m��Н��>�{��Q¯��FK����-��x����D~��20(/ ���<�6��.�U��2�����-�C�j���/p�����b|�橪|:X~�^%�B
ִ>[\<jHsC�a+0�dG�st�"�;��C��J�W7v��f"5�J �;ؘ�ݡVΟϗ�&�6�J���樈=���(������k��#HdOD@g�E\�3�"�MBR�!��P���B`�	9��3d�({O8k��=�*U���N�1Q4�bR�q�f{ݴ�Zo���N�E~��R��~�?3v�����bn�\#��s�c%H{���i,UK�nK�RGqY��y��mK�����&@~�_��o��M�	\������U���E&c�B�Z4��t�0P�x�FHv4"���3����#��"��{��¿�ʰ�D�糇��pͺ6��`�)5g�c�ׄ�㌌&�qt�vݝ�]jO�#-<x{�*>R͙���4D���O/*��4��b��\��/��(?��>R�
Ieܾ�#���\�M��	UH����v�nm][F�̊��XƨyM��+�$l��|����d�M��_�ܤH��v