��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸�Σ�HڂͨgT�W�1�.�gW(�CpzQx�E�.��4W��V���K)�����;E��#�� .��Ő;�^S�̤�WJ�b�]]>�C��i��¿x�D�G��US�t�::���ҫ��z	�p1�~���)���G��l�Jk�cK���Q��z�g���Np��лj�-P�e��H!֜)]>֫'����j��#��s�� Orl{��g"_Y��S>�E��Vs��_�e+B�_�yF�l:1BS���SY?�DӶͿ�(����z�\wQǊ��G���N����>��}�ܰ:��RO��F��f�>���)UEr�P �[��+�A,'�O`ޤZГ��f��f�%H�|�����e��yh)q�����ǇK i�nĸP-����"��e⛍Lm��[m�����T5�S��ք�)\�,9n�ޥ��e���[*�rRBC�'�����b����&PD<���7[*���)�����}���)�}�bM���f�l�:jA���"�E�pF1��C����;�9_�T��z*��<j���63��d��GR����?���۝8�՘2>~K�AnV��r5����y��)]��oqHd�=�6��u��}n�P���4F���W7�̆�	�4��F���\WfA��ht��d�4�LR`�	���&-�P%��A�s�Y&O�$ڒ�T�V_Z� o��r�9|��!�� p�T/�Փ%̌7�X�ծ�K)ta7�V�Ԕ��'��}��OC���v� ����ۙD�	/n�@�3tZ��4�T�zc�Gk�R% �G�z˦u���`m�$��,�����G9 T|����4��ؠHZ:pdW��!��X�\h�o�Շ�B��K���kp!��� �/>�<'�gM�؜��u�0꣒�t(�c��֒U����/��z�A~���HA{��V��c����Y�[4��'���2>�q����I	}�Ş�:|��Gw�����+ⲝ�Rۺ�NdCL�HX��_E�r==���H�"v��q'�β����f�ۿ"�B�r�ҳ�ma8�G��_(�U�Lw5m\Dy�	*3�J�.l=K����v�l��M�O_ �x��(5ad���4U�mP��z���q����<~�L�yXx�� �����"�7O3�!�J�P���uA�P��9R
�����fl����8�U{3�����B	fG.'�k�t�c E|Wo�s��gp[����4�2�ӹ|�N':��4Chl|��� ���#�Y܀:�j��X��պ-z̀D��������8E��	�!LK:yP�5UO���[�V�\�Ķo��A�ׂ��i���y�&M쎑��*�f��/�����.��쾪Rh8Ӛh�ֽ�����O�i�z*!�}<����XAd���`��j���	r�|.��C�n�7�֓6�ٹ��;�x�y�