��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���q�����W�E�9 Vοօ�̷�S�;(B�����",�U�s����6���i	t̂9։l��cE���	����a����	YD����g>���\GwB^pI�wż����hP���j!�(ص0&Q�m�`��(�Hd�j�Wjc�l�s��Z��^�V%���mT�,��m�q��a������mi8��u����iR�U9c*�ܐW���C��<�s�t�O"ˢ����m���KJ鸒0t��O�2�Z#����\kY���V�1ԅQ�@��w4��48��yhiz|+�Ӷ�r~A��r�MV1*����4����6,���Q� ��,�ܰ?
]�uv����|5�-T����DD��362�U��Rmep���ѽE���C.H\3�#h�ٶ� ����bþ����Π٣��UOn�U��y�- ���w�a�T�u��`Eh�$(����n6����~�pU�\��k��RDr(n�p���_���t��b&Ċ��-9ޒ�a&�(��z�B;Em���Z���9�r��d��(M2��r{�v�O,6hU1"&��_I�I��|��-{;��t��W]/$�h&�h, �+d�/�H�nng�b��e�c��j�5��m8i�����{�ު፤(�
h�����~ ��m�����e=
��6�D�V&������M�IAin�����d1?��SB�$�7?vy��@N���A�2�[�CN [v-ia#���ձ�c M�ҙ��/l������Īk� m��Z�Vl�#���c ��pa�ӉJc	�RF�A�gxl]�|E��{5>��`ޡ��W�I�qwg�vǕ�<��D�*��]�5�����^8���j��j���o�Br�I"�y�ct��Vc���9d
�^_�W����r�87`�:V�50�Øj:fK�t��l�;�*�7�"�Ro���TZ(�A�y�<�F�4�/���pi�����Ds�֠$Tu��»����}D%=_O��p���og^ݡk�t�dX7z�����2����I�(�̮��ˉ����}���3�������w�@U.��6���$���bWBVkXd���a��b�%�I�70|�)p\� �L��h�?�Uj��i6�\���!x�8l������sQv��H7��4o��)q��v�N�}�E��o(���F�J�׮���t��/�ŕ�/���Y�ل��T�9�^����{u����E0(_8J'��� H:�0X�潴e}���I����\��/.mኪ�옞Q� ������S�kK+` U|��c�=A�,�/u��F�7>i}$HJ_�(,���ۨE �/�1S^�4D<�A�r���^�aObw$�d4s?iCN���(�����U��>�ĂX1Lg�:��C��t2Fo"
�4�QP��Mվ���ˌ�D�<�=�KL���_���E�[�A9Ļ�ʲ.��^I��I������b�*��_��&2S嵍���+-��^}W̓̄�vH�={a�c��7t��J�0My�5^�2�(����_��p������$^���K}�ev������QBƪ��[+Kw�l?��C���u|�p�1J?X�n��*��\�c��(��S'}������F���c{�."�Q�a5��ٲ<����
"L�<�z�Ë����P�N:�v��1;�ƽ'	QZ�ϱ �Uj��mՅj�%�Zm�����ǀ��&���c�L}���u�'���rM�)��UY�W��=��j�\h$}n�U&O�Ӧ��y����O�I�� �xC�/�jO.� ��E
������!��W���b�=�Hm�w>���Y��D���|B鞦�%r����d	�;�C=��f��$s5�gU�ˠ!�^�b1����C�Vjq�qf��Ħ�ܢ\��ͩ�l�Ov1��q�*�e���w1��>V�Ex���e?}����HHk��U����)�����x):��H����������禭P?/-CK�rP"ay��~�P�YC�_3�mX�s��9�s����6׫s����)���}"3ʖk�a���V*��&Z��m@4e�O�����s�����}\Īaϊ	0�n>ݹ���si�x�!�$�����*�w�͠�4-��%��5J��؞x�2YFo.���c����b!y5d��bc5�.�j��C]<aZe:��D���b��$rW"����d��U���f�u@�J��?�J�s��S��E��0��$�*�����UXeɸ��(@�Y��iX�mِ�o1Ղ���"&\���:�JN�+��h�W�?��W�����oΫ��&�6-� |n�D �Y��؅.8[Ҳ����ȕ�4CBe+]�z�B%�����-��^+N*ƃ���ԑ�8��j��g���'�J4!PT��J�(PP�DL�t�dc��l���B��^L���S��)�%�^�9����|>-׬u&"q������:@�|�����gHρ��C(�.�p�����#T��pQ q�zݑ*���_���T@.}��y�5$��_�Ƀ��q��}�m3��T��g����c�V�_�!�9�^j�S#V��l�:������!�����i���=�[v�YN�q w��%aa�[Ùə��b?js�j��11�C.����4�4�g7~��M�����
c�Tk���j���̶����U@\��U���aDq�ϙ��v�J>��i;����A�.��1� ����ӂS!M8�ۺ��4���XL�:������Jak�� F_<���LBC�%��U�mӼ�g�a%G�{�&G�v91
�Yz"�s��j4�m�<�齾^c�g����T|J�i��O����L�ٸ���d�6����}�"dH]�ǆN�ִ<?�l�U� ��iM��\��#~k�(y�$�@��pa<e5�Q���[I:9�"��ɦMN�h0����S,�񶲟o�	�\Xe��`Xӯn�*�O2!N�r+|w����$�S\,r�!R}h9��-҃�?��~�Nq�����5�T���w�/[���&�>7��k#$����'ξ�@Z�D5�
�ou3��Y�МP_��MgBPf3wgD��R
�/�Fc�)2� pF�ʭ��36�9�2W�$���/��6�*�ט�(`��n������in~���9�H�Z��gJ���%�f�ZJ\��Z#x�	�_�"|/�\�V�T+��S6��p�⯩?QOƱ���ܪ�Pt۩�6�o��9���K���v����!�yN8����q)F4�$���2�IO|Hb�d�t?�6x�U����b���`��v���%�G9%�pO�%�o���g����!����z!���U)LT����72�C����ܷI��嚾W�L�Ѝ�w�f��E�p��k��QO�I5�	rm��٦4��d��{\*��-��������0HNh�|���Q�"��	�C�`�YS��H�f����{���S��|m���d���~����=�
��v'�^v_���S<��g"x��A��)�Q<�*4�ϗ9�92 �ĉ�A?��+16��qq����b�SD��d+ܭ�V�)Y4p;������9��#n��+mx�Q�Z�0=�J����ۨn�ټ��;��x��,�LG����>c�>��ݦ�5!pl�C��� �dȲ�Ҹ�� /�igb#�/g,ML�u����I�l����d@��J��,��у(���p������/g�|.Kr�i��g&�F���RŶm���֜Zj���"Hts��>S*�g� .�nK��kݴ� G��u��'����\�{F���,K�{�ȭ�ˡt��ڕd:�5�,�UC�_ٺG�hx,tv��Jzd�o�qϘ�@F���w���<�G�:���[��QRF���wM����=��ȷ��k�2�NSC��xs|�cYE�-�l���s��{I���6f>�\XK_+���JA)H�2P$�t9
�Ӕ��ܡL�kAkbc�?YZ~䴁#�ѦY��q�EB�9�^�5��a]�-y���Vł"�l��O�^+)��� ������m'�6�{�M)��"t #�`sM��4퀁��3A�oΚ�p�w!���hz8��*�{3����ٲ����*Uqg�XWr(��יդjî�����cΰ�o�DBΚ�tF������3�V�w{�EnH1��n3��}�;����;yga��Kp��I`��u$��\�^��G$��/\���!�������>�;/���!�v0��`��׺�?,�~R���H{�}d>��������L$=M�Ë�z��\)�L�?O�����
J´���;P��]��˷EP�;ct���7w���m4׏�:ՐEC���Kt����;��J���&!�P'*�<5�S`�������5��/���.�\�A�o.�0�Ǩ�c�+�q�"}�Y������A���̨�10�r&��RDt���WEu��7��#R���i�1j�SY=��������W0���ʝ�W+\�{,�K��a�_�'^?#o
w�0��@O�_���Z��}A_Z�t��3g�s/6TG=�����7JH�xj�It
)�0&?Lla��xȁ�7{�?PKQ�3��61���JC��Gn �Λ���te'zO�;��6�5hd�cY�A<'�e[��~�W} �&�X�Y�u?p�� *�Nvd���I����W�� � �N|j:�~�EjMe`U������/�����Ƌ��<2O6��-#$�&1Ϙ�*����y�u���4�Õy�r��1��9�vS���p(��˓�-S,1L1��YOXL����w
�*�+/w�5��8�ӎ6��@�3ڊ�Jb��|���u��c��&�WC\ {���u	:^/r�0GD�7؊3{N9��R�O58��T0B���M��@�7ګ�S��j����	�ɇ�6�F��
���x��#��
��� �IS� �,`C�F�#I�A��:�D"ծX�d��F8�$���Xp�.����KLm�d#~��|�����D�2m!��'�>���gz2���e�yhM���j_,��VC��V٦��!K6�����l�d��9�_��ջ-hUf�@���(��Y\��Ʊwd�Rۖ=u=	�a�w+ŮY���*������lQ+n<�� ���2Ӳ))����t�-��[�>��9�=b��x��Պ2e��?����O	N�lVkr��)�n�%i���"�yQ�EjM��1�T~���Ys��M��{پ����T#7xW�	�P,K�ǌ��S��v>����c�2����04��l��(�I�&j!�Ct�3%��{*�����D�h�F�����͵w��\��	�?�L���&�+Q�Z#�H�r���� 9��x���.����]���|8��糊�0�^\t�l��Ԝj��&hw .�-^s��﹎� j�~9������lN�2D���%������g�O��K�	J�ο5Lg���@��cbq D��QW&1-���V���D��%�&���U[h���J;�e�3>v�e6��G;����L��R��p<�����K�C�R����ƶ�"��>��9��&�j�}�f�*%�2�6��1�#���/��1�t'��D�_�����}2i�������R�o��y�í�(p���Ӻ�O�TbD��1���F�9Z1��5nnf�E���_ޡ���`+h��lx_�Os��TP|z��H�|���F���s�6���lBruW��p����[0�l��T�f���v�viP��fve�2���4p���9m[��JJ�7Q��842��#L[Pc����c���}y��j�~��i|S
�HR R�;z����9G�_�a��1�1��P[w^�x�7�����h�;y�Tu��+[4��D��a�*-|nI	|�[C����;O�HF;ӡ�sҵ!�1�\�D�u�1��y��e�r�.�o��	9C��>.F;��r�Q��W�)0@��_/)m~Kz���1��2X{wH ��,��a&�G�]�tP���a����M*���(�15i�Y9�{����$��R���.LH��H��<h�O���2�����\K����JD\��JLV3�:˲:���8��`��l�Utp����\[N����@��O�@�ri���6�J �S�|��{R-qO��706�Z]LJ|����5�7j��fD�aO�7"h��덥H����'k~�kN[FN�5�Hb\?�s�gY�2���EP&9ŀ������n3��X�%���7'����۫��J�[(�>l.�SS��9|���˰VԊV��ܑ�ѓv�o��u{��ŝfKm��<����g�)�.�����{e��Z��t��0C�s���X�}����,Q,�����$l���D�{�4C]$š�W�y���W�ࠢ����3=(#Csѓx/�q�������
g�hӝ����Jl���9]�`Qv��D���2/����|�dΠ��6������5��0�%�̝�������o�z���rAB=D�+��'��>��xG5�up�!���pZ~unZ�z=����-�;�Հ\�{팯�B�h�9K_Z��L�c�$h�!��vO�e�eC)�':�u���+7Tu��%<�V��5�]�}K�Q_��`�Xx���g�ǌ�e���ՠ�0��I����W3��pWm8�ֽ~:�.����fnYm�~"�<S�.��)�9���t�0��^�ibdE��降^˦e\�Z��1��#GFrtcF���O��\�%в�-��i(���S��_d>얅���V?n��Q��h�;�_1��zF�m�Pb{�l����xGq�G2�9�ne�N�U3fIV*�;H�]��w�GOS�L7l���]<�)���|8�;׆ ���1	28z�R�=�� ;)��ʸ��Z{� ϱޑ]QNR�w4����L��I�(��5f�-o5s�w�Iu�pq�WR�	F�c d"�h�>j@��Uۊ�{��g�!�*�y��ŗe���\s*��P��U��xE@�
��! ���CE���Y岓��G��u �Y��|F�8�#>���N��m�
�~�E�:ʳ`2��3H�G�q�WV�ZN^u�S�x��� �~�_Ʋ@)��G�kn�}��#�|?20��a�N�ߑ\��U�ݕ)S0��g�){�s�܊���\şY�#�˧����kJ���C֊�M�ĦE"�����	��˂V�`��?��/{3������a-��1QN>�q#0�_������Bcb�i����aT��4���І �
г�����g�I��|��2��c�����ʔoѣ�1AC{`��i=�>��T�U!�@�cU�ؕ`����,h����Dqz&:_58a�����ײ1U5�/i3�(y��U�/����@��"�Y&k	���}-"r�e��2�WƾV��ٹTT��V2l��,�+���T������^�qg�#�N�{�]�4-	�����,����ޠ��.Q�+�*�q��g��=a|�_�<=�f<vN⹠�
x��Tv�{�?�C���c4C}��x��'�c���&)��YHŵ�p�v�s��(#��J�)ɏ�K����_�!�y��ǐ�o魥b��'p����K�շp���OB��l���g2����S������Q��!��)���r�|c�BY�Ǐ�ŵ��"��)N�8���Dw9�~����~��材lz�00��1�5��޸�u%�S2�H�_�'F����*uW���%O\ﱮ���]�'�O��I�Ś�9ַ��k�G�]�B�b�k���kuP-�.ʘ�_�2������$T�0��h>��O����G �&���|�[_��ǧ�.w� P����^<��6��������]f���3d�#(����0�RUt�꒔vnPT���79֊a�.8�uЛ6�N���٘��H�[�
�E�ܛ���X�_�r8@�yOstCCG��f�����+��?�C#bh�t
�y�e�6�!O��'9��L�vT�G�0��"=�y.�����M�5��>���w��[E�����ܝi�1����zK��;T��Ɖ��I[n��y��|�ُ�����{rj� ����^߾��k�	?� ���tЙ����	yI{n����R���ۿ?8`D���%���t"�-��U���z��fˉ�l^���ʎ뒾N��$�O[PR����f�{�B�XAN�|��&���^�y��G�ϩ�`,�P����'����h�"������z�-)F�g1q�t��cV�	hm�L�Q�8S���/�%�Q
��rPU�ֱ��f%9H�R����S�Ѫ|и���<�l�`m�l��������5 ��_�r%�#��3�#8�5�#{���2AjY��d�	Hk�)L<}�@n���)��tz�m7g�BxA��3j�����הDz�>����o� ��I�