��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸�Σ�HڂͨgT�W�1�.�gW(�CpzQx�E�.�@�6��"o�0_d�h(d�����lP��g�����zТ��Thw�	�1�$杁���8Etp�M��Fj�"�v�S'�v���e��>�2a�����\�/O�e$���A��o/C�$.����G0�c�Uj
b���RT0��B=��ʰI�N��d����Ν�R�y���;eym��T�v�@.���A,O�[��N�kUu��(lFz=�vAw��T�fڶSq}��1C6�����j��a_���ih����oT� A��������)~4�QTv)+�"z!iM#{�~Z�ê�+0��I)�{�Kp�������S��[3/<繳K	��M�7؉�Jw�n>�R`L�*s����E����8c��s�Y5���+��2�V�l;�g��h79_����Nm��j-��e�SR�|�����58�x�����q�`���^�gܵ鯎�1�/uI�:�h"T�dz�eeP�kW"_�]R�.FO!�ͭzdA!���* "-@
2
��P�Tk��*IMgW��|Gs��#1�i���W9�+C:ֲ�Z�B��V�Vkv���[��	�oS�,��ί�z@*����p����-�∫��W>����+	�-�kMo������[~ 1D�����W�-�K��$�Z�����$v�ސ62	����ai��)]N������G��1��L�(bQN9��B��J�m�c�!�"(����q!;A�js�i�A�F(�|��+�6݋��G