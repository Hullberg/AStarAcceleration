��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���qm,e9��Աuű���z�B׷��!����c�FӁ�����`������F�;S}�a�(��{4�4��us;`dӷ�i\�iB��[��X(��\���>3��C���b:A�U��n�<4�MD4|���wL}�2��5��F&D>-z5·ޚ��)�u�{�����C��/��X�i��x�� ��]PB�L{��s�-���uu4fyr��vÇPwz\��T�d�%[�T��}e��jɼ��z̾��Ʋ���o��Z�yYG�p6\M�V�<%��[!E��wR�� ��w�2\���N��;b�:�����Si�>�+�b9������h�2ی���d�aK aY����M�(���[��(2��2UaVἵ��c���3�rIa�B�¯���,�����!�}a��TC�d7��'*�s���as��P��^Z��T����gL��`Y~5�`��No���y=Zn�R���u\�C��Z�- _ ��o�j"w�/O�ho��˹��I]#�>���'[��ƔN ɘ�T����jC�g@�Zy
�b@���ts5M�����Z�A�'C����1�����X�_��wuJ~�@`���%xTne������������ɯ?{,.�9��p�遇����B<�QM/�Y���p\����B��9��tb��vW=E�Y_�E�=lx��,�F����r��K%iGb[|������[��n����>ȟ'?9����~��n�W�ĀA���H%Jt�JE��б?dR���Y{^m�:<��$z�p�%B�4]wB�w��4kP����>����ߚ���CAω�;G��29"�	=��({����@��H�q#	�1���"��'idU�p�LsM��]7	x:4���z�o�/j������___��$0�*�N����Wݶf��k.��8tl��U"7� �;K�`I�4�lO�Ψ�
k���KүՂ87�!����c<5��޺�s��F�X4��I<�B�c}�B����gP�M���.7�Y��;�&�2�0:��[�j
����� ��rq�RѾ�?���M�8�+�Q���L	�it2A�\��oOR�#�7�+Y��}n���gΎ���B���wu=l�A,��B���,��1}I��3�	ܸ���Yl�d��\��Mx��=&���7]�H0��o����9W��K�>oRd�ǔt{$�GZ�����%�����va,�C�����xQ�%�&8L�RΩ*��҅L2����C�"�f���R`
�2$�}����.W�A"O�������xy&���o2W�c�P�"-�6W�bT.���(��8M������ G������%���g3����D���pư+��R�A3#p|�<6r'�֐]�T��e���$�7a���[]Z�P��J71��2{__�y��ٔƶ7 8Bl`b���Ou�P��VY�{�q�-�Ŭd�g����:�����Io"��eI�W�^�� ��b����<�9�\�e�:����g͕X/��d�-Ab�=Ӂ�����X���Y `�c���q��U�#@r�U:��^-[�Q<�":v�5B�}���!"&��i�1($?�I�?�e`*��fǗ[����"��F��-��G-�'�j��hHh0<GNt�Fq���Hդ��9{"��w�c1p�����ǜ����1�^����}��q$��5��}.�}�j�s�'����fHx��= ��҅z���E�PR����`@��&谤�7#X4��s;+ry���1���1ƶ�g��dOwU&�,0��;"�ˁi{ov �s":��Eu��R�w�Ij/�������V���ͣ�AH��Vh7�.�UOm�4s�5P��c��|���ݚ��}�z�l
�]~uFC"�)��}���J��Ul�Q�,<4K���dt������pi
��|��t�Vc��}��Vc����8#Pg5���3{� Ձ�Jj����2�b:ɶ�;[��[�KIa��k��4�5�k�:�,��>;����?�t/n�[�������z Jx�
��gл�RCg; d����l[t���m�8í��*0�/i��&�� k&§�C�l�,����~x����}�Y����Kx`&��0[�}w�:5|�"��Z;9����j�"�K�l����N���M�׫a(����T�����w��]�𝝖�f�����"8��E��*p���lDD��s������zQ�݇ݍ�qA������y���