��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���q�����W�E�9 Vοօ�̷�S�;(B�����",�U�s����6���i	t̂9։l��cE���	����a����	YD��x$3l�k���HWs(a�t��v���ɺÙ;t��pl�I���X�t ̦J�����c�0����4�k�l�dY˙l��!i�������>b�n!�+뇚i�=N�Y�,���bT�zD}�%ߌÆ�W0Ǻ��lw�g<R|��k%ET�����%�T��9�s'��CX��~�(q���� �X`ă�t�C��Q؊�g^�s�O�}F	���j�O'��3+Q�*Иt�o�y?��-T�;[�����'���Q0��@_�����]�/�����~K6j/��o74e����~ENQӄ��(E��we>m]]kU������O�A���Gjy��2۽��V=!d>j#a�q�H�sKe�g�^���c�nާ�O�?P�zo~� kARD�{�-H���Se�F��(ZMT��D
Ӎ��c4�3��@,�,�O]�g>���.��KJ=~��_��z�xxRG���f�u��y5�p�E��.q��	8t_�q5B�M�p�lK����3Zr��^�������#"�9W@��B�[���K�U��ٵv��!Β�D��	r}�}J�n�@iF��ӧg@O����\��{�
e|k��`�=��\6%���cn9������W���/e/��+BO ��_`ǳ?�+�a����,�T�� �-Bf�d�)��	O�$�#�X�Q&c��l���G�=�Q0��DP�=���Wf}?tG����R�f�����k�ys�q����np8�IB&N�~��tXhO�qǪ\H�T�a3�V�R�8�;K�Yu!c�V~���}��9�+ =��Rz�k�S���Ka��4NY�J�,���J����1�I�������xO���(Q�,�O�HXsR���.{D%!��~_��{brJ�q�����*»��W�ҳ�@���q�=�y�	N����<�TUQ�}�E*4���j�Α����*}�j�K�ʉ� u���yucg,����C�uw��}��8�Uc���3�L�ǳ�B��c�.��,�Ӿ�����P�9)Yc�Nu��?���j`�U�d~�?(�~%���/���Q���h�d+G��!�e8��\��.��B����A���բ��%s�nOp�����js�$��ڣ�B�'<�k�/3o��Q8S��"���������'�}V�6��BfQ����Y��WPi�)\G��@Ļ`j���C�.�Z^O��.��3��]+z�e||���Yq��FΪ��M�3�U�/=�{��">&ɏ�� ���J�a]Q�Բ�Od�4h��:�
�K�.�0|lfġ�_W�CTd�;Ch,JΟ��G������}\ ����L�}��j����Y�d1 x4*4��:�n���%�%�VN�j�gOf������u�b�{�ܺj���h"�j�K���q��Y��Ő1�Tl|W�����Ƚ�*���8<����7�!6[O�]���|u@��X���Rڼ��+o��AU�6�6���ccwA�ϑM0V��x������L5��W�x���5�-�6�������![&W�gv�˽��2=��.PQ�)��`*��ao���W� �G��^;
og7���	����+��ݭF�_@���u%>�E���t6��;���p�[�(��s)0'��!�!mz������Oƅ\�j��LWp����>o�M݈�˅�W~k�$r�lQ=�/𾧚�W��̩|����k6+� 4��_��7R���H^.X��[�Z\1���Io=��nj�^�LCg\.nW�i��9��rM�'�ig��)�E���?�6���X��,�]��!0�$3���e�؄Au�W�hA=i$��]���J`���v��gc*�D�8c�1Z�J
�Z#��h�_��(q�ZB2�K�#��7�o��-�o�Ͷ�uJK��X�$r|���f�Xp�+�8A1W�Z��0	1��x�[�li��k��s0pY3�4�N����(¦3-Z�WsC��3y�V*k#��pQ��cX�ߞ���N�	GT#3���r�(��
�ԣX��Wʈ��N���6�o���F;낄�ϕ��b=��e��?����Sr.G�*:e�s� ��I{�,r^�C�iIk!E=-/^|�����G�	��ƥЗ챸P��)��[\���]�
ƨ(F�S7��R\I�(��R�h�q�D
�I�׍5$��Sn�B��������E�_��̄��x���V}���.��~�#m��4�9�i�N��f�(����"N#�b0�%���RR�-*�߃����3K�##��*$��11{{j��q�t�y�,�q{_>DS����1`8TY���#ęg�OYɢf����i�d84:��0�8&W���2���dXsemF����#b�Ұ2$L�[!���>Gw�����x�#�Y��Ô<���՛N�jp���˾=��ؔ�:H�WB����5A�X�?����R�)H����ٓTum�	{�Ԟ�������OZh�&}q �P9�������</d���b�/m�(<_^M� w�m����N�3b���>)�&�i�}
�?�Qu�0=����KԵ1>8�]�h\�� ���HgT�RBE:ěnlqD"%����V�8��A��� e�!Ҏ�|h��hZ�ݲ�r�0� ���L��_�N�v�c[��~#����7f�2"`��:߇o�ۢ��cU{<�昚�~e�C�R�@�k/������Uޤ��}]�����b-��	2$�<�V	E[1̡��9k��܇�W^K߭�e�yn�0iX���bn��������f5�To��z�ye�d�M�k=�m����h���mW�4��A.9Vq�Ly(� �[����,��M`M�EJ��_�����@��]R��ɋ���3X�]����?,5�N���0(݌�xL��nX�W_�]y���H�]�� �n!��}��{���he�aaY+FС���>k���Z���IB���w��:�*�5��%#�����*�x� ��b�|�%�Uh�m�4��OUr�7�E�V8�:H?b+D�����7Y��qj�5���?\Sz#nCg���S��u��5��1��0�9��^����E����sL6�͢�G�����<K%���ʉ�>���7 �8�q�Cg���:��ƍ�����ʻǏ��ܹ�7m�TI���`y��9W�/��OL� ��i�f���������q�6m�ה���aI��S���Hi,�)!��m��WׂH���'&�A��m9���쪳���,ަ,��(�hzn��b�b��o�-�B����I<�.���޹�	�Tl��@9X�υV�����"�M�h�[�|$ئ�f�Rk��\�<q��R6�[�+�H��Lj�5	0N8�7���/j���]G�d�h����V)���^|�#�!W7�'��(�{?Y����=�S�W�t8��刾���#�Yزë��S:P)����~�gf����O�ܙ���ӓ�؁���+��J��g�r��׹�ډ�y��t+�ѓ���/?�A�G,�R���f&\]��{:�*wE�L9������`�=���c�뫭�s�z�����,��Y%f�T.�����Oz��]�>�����>XI�H����A	�Tid��x�R��FY���(�ŕ�K
q�A	(�R�!�סE=�@;8:w~��'���h�x�s���u��}1��%!#��&ř�"Hcs��~0�4fӹ2�!LI��Z>���:}n<� ���4SA�	��,	�ĿY��bk.�^�O_rM�K��WW���hkK����M�l���oE~/���6�G����-%���9~��l��^P˔;���'娵j�wsZ�4tJ�H$�/H�ZE�q������pC���8��<�����k���ic��om%�CgJ ��M�`��D�7q�$��6U���]�/y��c���	�D�!Π�[5"0���{t�gF���8����C�А�Z�2�Z.�:��~Tv��W I!���+���
��}���R�y���^���k`ǌ����}��P�T�0߄:�