��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!��ߌ�6�u��S�`T
��E�E� -�5x8�ym�7�4�����Ƹ˲[�B�?�O�a4�����ȅ~��>����8.�NSTiӸ-s�M��(��'�Xh �ܾ l�Lz�}�wb��=}�5k�>�b���!���E˴�O��"��ߒ�?�I X�"R� p3��*���l�.��}`�˷e�	�ݼ��{S=winDO��N��́+�����W�-0l[�k"�-+�Z�W��Z�?O�(&�oR$�����?�w?^6-�����0�d�%='��]5����#���͉*Mvb�hIu7�����ක[G��*&-��ݧKs�ah��Z� /��÷'j��C* 3v��a�0#��>�	A�������"�����v:��n����H��BXg��~n�]YRK�D�y�VmD}2���@MP���p�(r_L��W$��b[`B���d��p]&�=��H~�V�m9Ц@!]��S����T������T��π)C��9n���rĐ&�c9��'9����*3f�!��'?܂�������͸^���|:�>;;�Q��{�&v�@4����Ǔ�1ЧW��I���*,TP�/@����2��t�(� T�sf��<�����.�k�8&�m�6�d`�eU&����Z����:��>������c+Q��eu��v4�����u���y_�c��)��2��<�U��f�Hɞ&�q���	�,�_��*�XA��O*�Q�O�4[NT����}ld��c�<+����v��a�\��*��^��n�������}H����e�T s �b���d�\_�ƨ;�W�¹�?��yc�b��Յ���<��6!��>͚�6��6����@�C��v�M�A"�=80�H�\��0�Z*���O�a �qzI#�[Oӥ�LO���l/���Dt6�a��&����>�������Drsd�A��&)]���c�a����]�6�q����u0�������e���z)��n�cl���0)��>��%S���ڿ�b���@���ky)R����%0Ŗ��`���#����λ�­*�	?�:���\�����#>�Q��:��1�?H��2�C幱§'{n ��BC���Z���'��2e��Y,5C��YR)��0}5�M������ߞ$@�r{���ܶ?_�T>bL.�=�Z�A��~�J�{B�<h�����\C�M�m�1��i�����c���OW��e;2��ӚT�t��>��y����-S"�����e@X�ch�S>�+���7:�B�Ɏ]��A�k�<���D��A ��9���	 ¶�s�R���v��W&	�M�M�23��G�k�55L�[�*���J�"X��M9��y	�$y�f_8���ڙ�SKѯ�3����F��Zؤ7 �$#�*��Rv�P�w���dCۊC��i|D�`kZ78������.M��/h���zu'V,4x����?Х��{���Y�	����0��m��u�~�R�	�()��Y]N�фSRGs��y��kK)�> ���HS|��� v�4���!��a��RI�a�<r�s^�X�(�С��\�qcZ��$U	�� �&�=Ö��?s�a��=�f��pF8�-[u�ҭ�@@�}<���o�����}?ܝ�;�Zi�*�S��9��<����!�WgD]Om���;B��`-�4�.���'6��_L���[â�A|��XZXd�&�-Y��,Z�J��FŖ@j���^'����ds���nU����:&�@��dʯ8��2�$3եd��*�U�-��0�svT�١p�	���+m��$>&���oظJ��M��P�-�����܄�f���H�T��S�3��闠�h��œ!��'w*���}�X�&?z�M'�\T +̲��Z�.�c�m�@M�RZ�G��tk8=^���ڀ�9G�z�hh�7�x{��b��e*-���ϋ��N�����~;S,u��"�}�;������G�J���߈�o�Qh�����?�̱�c�ݙ���$E�B�x.���~-�g䆰@�� ���y&��	;g�J<�p�,���Ϙ	3r�g�I��ϴ��ŀh��IH3��#��y���ul�IG���L��kXӼZN4�;6�������TO��@�^^��a�8�R,u�޻�w�g�vP���r�%�#<�Ӎ#-��cj������[�)>��ϭzA�ғ�=�n%��u�z�s{��NvB)���u�Q&0܈��5@j��EL�H�h�+#~�)��LX������3ޚCc��v16��B�I�}8���V�;S�[+��N�f�Ёj$52I��~%�"�����PJ��j\���#���b`�_rc�ܰ��Mw�F�|��.Lc ����KH����nsU�<���e�C,uJ�a8�va7���e��k��
�{��xA;��D5BۋJ�B�T��i��H�q�=ˊ�8��i�\�u���\��9]��K�j"ږ�6Z*Y@ ����btx�L�_����\4���eب"iA���E��i��K��i-��L,��_���8h�X7��j�Wb2�f��1����͒C2'���p�B�ɣ���%w]����2����ҟ�*H�Δ�+n�ǎcx�̵Ȋݨ:	?=��b7���<C�]��P�Ǩ���d��bh>r�];v��\�ɝצ�&�����&UtL��z=x��E��E���R%87fb����ӻ)W�\��wӶ.�~ߙiF��U��P6�q����%δ��<t����g)h.&��N@r���4#��}Ϙ�rj�0�?��K0'Kv�5���.\�.����5f����J�rd�B�ﴞ�Y,=/C�X)��d�'����$�J����<�{��V��8cĥ�j>�����^�q~Q�&迊���O�Uc�#����	j���tU�d)y���$VO�{�/&:��@��q�����+�SeMc����
��S��̒�ɖn��x�0M���W
����wР�m�2���k�M���Ã���%�b����W���R���q���n���cZ:&�� ?��Mu�d��W���㸖Xˠ��k�7ߛ˱C�p��j���]��X��Aa�E)��U�,���*�s��;�.w3~�� �/��P�݄�u*��#]۠9A$��ԝ=��S�k��n�5�AQ�N�W����]�tw�HK�3�n��:M�ׯ;�#q'�ЙFޱ������dk��?��X2{��2g�C.,���<��D-j$2*���(�,}�q-�TD�U��'��.�����b���{���ȵ��h���].lh�(�����p��� �8��M�nhؔn")�S���_�fdjZ7��J ���ePF]�U���h�i>�B}����0�N}Y}��}ErL�˭k�oUS����w��ITM)"W%e�)��Qw�$Ȩ���l��x.g�����#�6��lM۟�J木�����*��C�kS�=a�k\�Ɔ\���%�8�������uI����hX���	r!֛L��N��.q��X����*��1W���]3E�?L`J�,~Ў"S� �H=6���Qϋޜ	 �0@�r�F�O��P�,��������Pq6t!�Ґ���:m`h�q�q���wvk��#���ٗq��R3�ۺ��/D�ڟ.@-Πp�߸�u	�'0"���� K�N�����Y`1��F�.��3��E���f(oC�� fs����G�5c���ls�>�Ø�*+��#|���yUi�$4��!��~]��*|e��L5!����i��Teg;u=A=P����M��"�k�b�ϟ$��u��,�?Uf$6�Md��^�"�I@�FV��ߟe�T�(DB��S���f��V4�[4Cٟ0R\�.	� I��J��,׮�ݻ��g��4�#
�?�*��me��=�2�����@�S�]��H��Di��BVH�b���Ph�ř?��`��1��� 
YX�ALb����LC04M|O�Ԗ�f_� ʤP����A�H<q?��='�|ts~�z���M�a,]��6�(c��M٤a�\%�iU�4R|�^�'/1�ѡF4X��J�$&I_loؿT����%S�Q��߅䉘�i-���^`��64��)�hb-�r�ؚi�ʮU�}��O���9J�����q
���S�p��+����GY�����/F����Iщ������b��@T�X�x�M'�:�k�L���9��!��Ry�����;��]4�D<�#�[��v�+�<��yV޿���1ҟ���#\,B�V��K�jҿu"A�<�L���kь�~�kZ���s����M�j�B�i�a�Ъam��#҃�B����c��z;%�õ�o�od�e���"����d��.?����5�Y����u�*|��M��hV�- �;"�mMk4��ғ�X����.k����$�2��(��1XpRNeS�h����M��͂�ʟ�F{&3�>�n����?;�'�G�w� Q���E�@{5��%#�th��J֗ �A�'Uq����|f)`Ra�=�´��ݼA��h�II3�E8��A-���HE���Ok[<s?:��DO�� ' ��;X��e��
����afa�A��Y9{�*08�4�	.fA\��Bn	�<����,d���
{�U������ә�0�gd�&�-�ń��*�na��Ԇ�9ׇ�0�H��s�ů%���$
���)�~b�=�U7���U8؉��}#c��h�?L���C?xmg��p7-��v��L5���͝u�I�9��ѕ�@h�\%pc>,|t���a%5��FnLU[}&�����Rl1����Ƴ�(�{n>fD����ѡ<��y�V�ʗG8G1��:�	�sܻo�P������l��K��N�o�kKp�q'l\�k�5�Mݭ��C%p���|�c4辘.��Dp�]AC@�X�۷p�vh.���D�`J�Ӈ۶<AI���u����x���/�qFl�� �Ytw�dK�W�.��dy*/�o�q{��O�K=�g����o�l�6���6qy*�cUŘ�x�́�Wr����q?P��� ��o%���.����(�,VГaf�h4'�^��T0��v/\].8!$����me��K�5���T���M>`�1��'����xy9n��@�}�q9�G��ҩw�AĠ���q��.I��R^��O��������V���`���4Q6�i׼Ar�!_������=e'vE��X?607j��.�KZ�1!�$��%m��$�s}��n��Vx������=�,�B�0H#�~L�JT�
��MD�׍�Uk��p��,�����6�q�W�25~�˫s�����P9��no	r*M�&*�r3O�3*f�]B�y�K_0����4��� cs87>�&;�Gk��l�/_�H����2Tv[�\̼9_Q��
I�羔�:��nKLQ#�Ew��<m��U��|(���
N�O{���.t��E�F*Z��'#Q���/jA�ڌ����@@���5�x���{"�B��&C�^���k,U�� �z��"�=[��sD���+�5E��,@f?/�J�9���������/acr��o�ʉ,[�`P4^�H���ts4-�e��:� �}Ja0Ō<0��+�DQ��d2��<�;���܇=�$NC�4� �O�!������	��\+Ǹ�1�]&��d�����:�D�MU:*间W�M��W�*�Q>f"V�z��*L�LbVWw���sYR����g��< t9G2��U�,Ұ�0Ư�kաBAp%E|?���7]�R�G����//i2��#j�if��܃���QP̡��+���h�sW)*Y����þ^�[MO�-NE�fڱ�QՊ5�Q�xց�G�"N�$��NQ���9׹���~��I�(@�۰L(li�?ē��-���gU�����e+/Z���G'���E�����J*���fN�B��������W���j����.�h��K����}w�b��)�ǝle�9D�Z۠���`4D1�7��ee���������4(P3�ԉ^��!���<ad����^�.����W,�C�D��QV�]�`�̉����֩�ay ��"p���[���,$�sl���41y5�d�Y1�cF�5����(݅��r�_�~&;��m�[ӛ&�-v�LYk�S-��16pß� (����9�؉���˷�N��j�V�����	'א�V���zK1y��)�����^��P|�k���p�UT}�Te$	���g�sr�{�3����S���3`	��-iMO��o-�=�ᅑ������H�rh�#� ��� kM�S���c\�Q�G5��y�CY�T�j�[W3�MqY��'̼�&z�ڈAfI�m����YC�mv��n4�"�"�w�W�I��& T,������F��a���DD$=�[1����`p$>���%Q��h4M�cl�1'3����q��>�m ٓ�܎/���)�D��wfs\�x�!i������g�I#��u{�J5���I�k�ڼו��i,$���r4S%D|��d�7���
��ٿҔ{y��J4
�k�L����.͉`(����9B̤��Lh�vw#�X�<7b���5s
^���c@�i��K�uc�|)x�~�%���6Z_�N9��	����	�n��a����R����.�2�7&x�Wy���!���Eo�7��K9��j��Vw1�qؚ�o�*�ׄ_��}�#���,��b7�} +:�����6�=b8�v>��C�Co���"
ގ��AIC�It��J��T=�;�?u�r��-s��9xu���o��ǯW�x�X��п��6�ϗ�P����x��̀h�ѶAx{Ȑ*R������6TY{J�׀�t�&�*�U��O:�߬ � ��B��{�~�Z�4^�-���kpWɹ�4�dw@����S�����>�@����$�y��*�<8�x5H�"�ܟ�yT� �q|A�]�D�����m�6:D�nC�O�	9Ku�D7����ˍ��o�����]5{kB^�-X|69끖%:B,�y�KĠ}�ټ�5J1OA��C��?����������0���� ����稺[���R����v���x䦱r	G�:Y(�$>:�Yғ�
z���+�y��%2Q��m�(#v<����Et�BL��w�8�K�	��9H��
oGtǹ�����4x�Z�B�������I�w�f�j��W"��4w���%j��>�cD7�G�X �@'�����`�ٽ��8[5���k��:��bA\��x�15`�Y����'�g֙�e"�3����R�7U�YUu�\�D��A���i�
��;mMoDh��}�-ƀi�5�#��}(k�:5[�X.#߄�� �"9�&��CD�f��=����/	��T�hG~w��NF.��n��c�G�2C��qC��N$���2�m{u��̻%d��s��Rp3)��j�;Z�ʳ���͚a �FE�a��	e�'��V Qf�sC2GQ���:+�ӽ����P'jt}w��*#�C�D����j��k�,�|ܵ�W�r=K)SՋL9S����vF�H˥��@f����l�M�%��ܘI̒�B�}]p�q�������	�h_ۋ̺�#q�A�<'r�lJ��03��B�dE.�\���p� qT�pe�~R��E����Z��.�����0s⛱�U�Y��Mko�*6��q���Ǥ��D'|h��9l}}�1=��cox%�������dh�X���=�!Xo�����M7r�'b���-h�q��i�	R���/X8��@�M4=U�����⬶���G	��,����J7�A��UՋz^-�e+[{��T�!2Dn�P8ɧ�#�=���aѿ	oC�[1�>��u歈��o+�o�?{��Gוֹ6�I�[�2�;��B��R��	\�>Y�~�إ�x��]�'6D��(�ҳ��e,���8���M��׃*o�T_[[^��k��b���׍��ʸ���*v�e�@�L����g]���e����gԃ�!��Ce���W-:lvL}���;%<��o܆q�!��&�;#Zz���緢�.,���.�vs�f�4w ��Sȥ������ ��G�N9k�/�h������H�zQҴEu�9e\<�k�˝�-����4G�`��\�C�SSW�A�ugI?�@���\�4li�.�����l�G<��𳪜�7�AwNs�?�x��QV���2#����V�C]�6��f(B�_;����+I�i��-��#�B?�WW�PL"	�K�]�#�u��3�d��Z�u��<Z���@-�=V!7d[�<�_�ZA�XO�"�CW��B�ˣ^�[:�&��dgH*a�>���l��Rp�h�6D�շ"L+X���c��b�n�[�N�0��
���2|�#?����z���ec݇`�D	�#t/�p�v�|��	��L�f;�V����|�}�C�y�Kg��OB���a�K���[���k��G不cԩM�ut����<U䟌��W�<�nG�T��[�g*t�*��*����*���׮.�^}f�v��7w��M�v��)i��b��,��"^f%�-l0o~Ȓ2=%;h� _Yٟ�iBD�ۘ�DX�F1���ZN��2��E�pu�Zj��zk2�{���b@JOi;�Q&hﮘ���x�j�����Gd�D�� zZ���a5>gA}avk	���}T,K�F\c�7�#%4�E��K�=��gl�X�ڡ�)��ɖ� #O��	o	�j�L�0��/*$_m�s��:���k����7P0Nd�?l��b3<�(��A�7G�h�YZ�c����+~�����>��A��s��eS�t�'�dFȊ��6+r\rt��cQ�4�U�ӻZ��ꈞ�N��4@)u�(qq.�h���xڃ�������� ��̽�ט5 ��ג�!`Y==x$��X�β7�i�P��׹�D#�|���`{��5\�n�w��Gu���x�����Q�M��t�k,�Z����._�oz���������lk�t=�M�DvX��p��KW�ӝ�M}>�i�9�v����h�R��p��F�课!<�Y�)ΰ4d��g�h�����P[>kڡ-3�խު�r��LK@$2���hvH �!2��>����3z�^t��\�w>��RJovT����45�E������-��,��� ߳�S��8R�}���}�M�S?��)����
��T�>�LB�|e�+�8��;�<�ݞ��^���v�u����JK
��رk�]�R�Y��z���a�����N7G��3��R��`H�~�2,��@�-�nP�d[5/:��tǌ�
����_
�-�����姕�*���aq��vdKD��m�k�}+V$T���q����4��|�x�y(Q/QNP䖄 �'T妜"�v��]x�c�M���}�`�,v���Ǧs��3=�������p쎡���(��=
?����)�n�SKH/�xxh1��Wk1��)���p|�`��5����L��ݤu741�������l�>�igp��0�Ԧ"�1�!��h
��"�Q2��@:��� _ހ�'��w���i�n��s�V	�f�꒩(~ۨnS��������n�K�^�8Rn�em��P�I/:���u������\�Y�П�3p��|H�KI�o�{_>CJ���^�5�eo2��}0�IgzVc~���{}oA��"0�2ޭ}ji�,7��<�U��.��#c��z��K:�$c�
��8��A�Ӹ�ɏ�Y�����h���y)_����qY�x�V�����g��8�+�3�+��oXPXӪ�[#N�T+��������Ԁ�J�B�!d<)�/}PӮ&��cgɂ�Z�u9gzA�mc��KS��2�,�Aޞl��Ua/��mgl�	V}�$|�-X��k���;�'� ����J1�}_-�v��"�@���@P2t�k�I�ȖE[�:�ϣ"�{�y��aj��h,�j��EƭW0�V5�Y���.�ͦ���|j����H@(�O��+Є�5�riJ�j�g=�= 0�"�h��s��:�����	��	������ެmZ�����' �s���pF�#����:�H�"|ܙT�R>����Iuz�p43�Ua ������Ih��q}`n�[�坓<�"m�q�8�¹N���ZNVʷ08���]_�hM~�loAy��}y��:�]�W�\`Ȉ{~WO�&1V? 2�.�]d6�J�����/)+�1���n3���-h��:n���X����\T�����e�v��3�nXu����n�X���˥c����#A�l����Wx��%����u�"������˛'��>Rq����DB����蚁�`/��9>��3�� Ћ�H����;��3	k
;����HNBmS�~<)i����S��|�L�����qI2��/�g�p�iL����\��&������D�h1~�N���Xf����l�cd�fmk�1륟
�y�iD%�<���_Pi�iN��C6���*z� ���6u+��Ƣ-�EEk�4�?(*�Bp���Iik�v�w5Eo^�I��:�$�s��0WB�C�sW���c"46Yح���C�7�纍���:F.�������y���O�ӤU""�ru���OR1��k�9��U |��J�~�+��`6�5Pq��#(_��Lj(��k+��s�z�s�{>���f�ܚ�x���ws��$
Ʀ)b�� �H�E���J�m���J[�'�hG҆i�\�`��ߐ.�9U!��T8�糅�Ɓ7%���0�m��Ƨ���73�qIF�f� �(��q�'Bsƕ���b��Y�ZN�:��"�7�i��aO$��!�-�Oʁ�>1�M jthů?�ϭ�V�����������h#X_���N8�9�h�by���l��v����g�v��ya$e��6eAi�ǖ�T����:=����J2���so�Е�.͇�s���D���&M߼V�Z�Ж$XL�ГF�~U�!4-��']4SYÕ�N�_Q<>N�w�kĞT�4��I��dL���f���kQ���څ�|'���B�2Yeoz��]`��5�ʦ��)�l�_��W꣺��o��ّ!"̼���H�Ժ�[���mh��Y���_a��}�(>Q!��3P�)K𩠝A��zc��㐩��x����[?̠����2y�PqI�Wq�
t#��3�a��<�ؗ�rNy���$�^�&��crtse�0��A�F H��F��H�s���'m��P�eѫd��Q�x�}º^�E��|�Vp�"y�N �eQ�'����n�l�¨� �3���T[�Uǵ{h�נ��FнK�~��t��9�h���ʝڣK�>3/�
%0�EڹZ��?�z��Y�Ni�R���]\�w��Ŋ�^���9!��#'����;�\%���ߕƣ6R�S�(��(���1�T�x�'�rϵ�� �ۓ�������ȷiɬ����Y��+�c���%�6��B���!�ͮuHu��g(��>u�ߝ�T�~[P��j�ޙs��$�����b�w&q/B�B��C�%��?��Ez�_�Q�Ce)6l ��Df�:>��%��I��7-%y�ﷸQ�:ZtJ�K�ݓ�s�k��D�}�u^�m Ӯ?rS�'~H��Z.6k(� ĺ���4�ms�FCʋ�o�&ڋ�voe!��9ņ�+Ǫ,���φeHc�2��K�}�\k�ѵ��m�����bĬWˇ'i��#�u��21�����\�2I�(�4!��Q<`�	�&:�_y!e�Dŧ9���]5Z�Sؗ-�1XN+a2I�s���.5>��]�D00TK��ys���2p���7C1��9f|��ZxuZ/�]�,�j暳WM �,R����R4̠-���.mw!�u�ÐNa�eN���E�l� ,�w�9 �v"=#���V�@I�GI��J�Rі�\/z�]���������gz�K�-���񕛎$���̋f2��nR�#�i�v��s$�X���:��!k����d]�-�|��S�hg��b�!�qs�����|ר���B#��Q�\���/�F<M�\�s(�  ���m���1 ΋�����oGA�Jz��(TN��Q��%�>a�
��q\a�ݛ�dDP��ץz�L�] &�,�я�>�U���������{��-Q�+��J,���`����
��Ca5�<�c ���?Ԣ�C`�(�!vR	O�Q�4.���-�B:4�uӖ+@�2��C��kP	�j��%����+�t�]����rT,E���ʹ�X�r�;ˬ�G� �5�B�T�=������5�2� c��+.���T������J�ܒ�|�B�Y�4-l����nK!�e��W`�~����Vl��D}�� ю԰�Z���$AT�2����K#�4��"%Xn��h��6��<��+S8d#:j`���<"�_�"o�L0���B����_�m��ש>>��b7��{�P�:}�����e�R��9��O����)���}�o�NЖ��xMF+�u���1���
����ĢPզ�MjkˏP;?��z� ��OY��zGHb���%�
�2^�s�
MO(~#|8���c6���2��X:M��A Z�m�:0��J��.�஄�v��s��+)�a�\��o����U*	��-#���A�a\s��-i����wA�uk>w�^�b��u�qXD5]j�nk=u'�o�݊6��~ih��%2L��F���z��0#_�����<��[��9����SLz��9Kk��^�)����7��1߳aC��Jh�fy�׿�b��u��Hܴ����/8��jtZ�P_����<7E!�I|�P�,Pjy	��~��:�<b�	���<n4��~�p���eT�[�4�2`@��`�g9�� �Σ��skѓ<�������ӲE�o��؞l���#�v�,��#��9�FАk�ԄZ<�}�^�\���C���ڥ@&�ۥT@ɀ���)3��44�e<8�P���ҡ�Lf�hf�k�d�E�S�G���YE��+^����ZSn�������J։�#@�$��cI�CU �Z�a�9��t;��e
��ID��{8��J^�Ck]�0�ȥٽ_z�Z�7��i��+����P�O�"lRoR yM3��|;�u�imwɌ�&��q���l�a�Z7*�e�s��JNP������j��Ѭ�B�)Q$T�s�6=�8iO�+ןゾ �HVu�F��.�@�=�u5)��xt�5䱻C�8���O_J�?Z�ϯh2��*/B��fl�|mǷ}�6�UnuhA�)��l�A���ѝ�$�ץQ=(Q�Ng�W�^���I�[���.�0HuZܲ�u���U�u��C�"���"����!u����d|"���vK�Z�fGf�	��1�ϭ㎯�:󾖃
I�%U�Q�||��Z�IE�k�����/�v���[uLH:Ɋ�p"��Ȕ5��V�+?�筸(��U����f��y�͎۰3��0K4�2�A)�n6(����k9��K�Z倇d���� k�7aA�&��j�9��'��2$1�c#7��r�s�ƘkÈ�~����h&�b(��I�t\�W��3�)!��A)�k�*
�\��!*���pFAk<�F�2�4GHe%Jΰrщ��
*>��VȐ(��joI��#Z�}�e��xi���� ��(q�B�G���|�͎L"�����t��oA�c��-#�o�f{��)�h��C1xW�9�z�;s���1���ʵ�@�Ń�m�*6�@��Ñ�j����j��>;���E�#��6�b=��0�w���XȻ�,�غ���G�*_��o�-)��%M �h���+g�s��I���pz�墊�!(��^�"�_r1���80y�>��SW�x���Ö-� ���W��}5����ϟY���}�gþd�����M� 7X��*�GZ�BC��@�@���w������-c]$�;"��wz��J{�	=X�-���B��Vdй�}\�=)�-%�eX؈�j��I�,UK������I�;h�������Z����h��l�h�N��Ƽ=�|���o�9�RяCr,��5��ω�]�L���14�Y��[7�1��i�4�\�w�iX�����<���$��iG�Ȅ�@���t,�E'�����\�`�d[pG���c�E8�ěNE �|��O�Z��=�;�����#�F�r��w@~�`��Qtkp�;�xX�����O��:�2g�s�U�s��Y���q0!IW޶z�/�� �R9���E�bl�{z\��,A\+�JG�щ'Çd_��A�Zw�s��sl��1b�����͡��e�=1"S���$�`� ��x��\8��"
#�|Et�����0�t�`x��i��^�l�!B�O����(�N^�CB����z�1T!���[��7���JjQŲ��ɍ|�Xs
�%��fh͏��V�c�.�}�J�p��D�\��޴�	��Dw�NU�Pg�p:�qeM�h-�0<��&]������ql��g�WH���͈��[#<��F���a;љ|M�!˗��t����8�����<�$G�r_����D�Y�k+��b�0�8Yz���ڮ�>�#Ī8+�^�ѪMAB�>���[�6p���Gc�e[t��:�2���`���2?��<�4	���_~={ S|�`���vJA�j&� ��=g��>��=b�H��S56��N���� �|�t#��0��q��^��� 3m���S�6��Rhw���A�S��SX�Q�K%�����rL8
\�c��I��F�[��ё>=_�6W�=�Vy��?����[_j\��^���*��36�a��D9�@�7_���A�k�O�$�У���u{淯���}�Į<��*���Ċ0�����@;�{IĔ͠�dͺ����~f�^]i��f7 �4TӠ��m�O��GJ1b�p�A����F�,�V���%�	:�%�'�Ƀ�B�0����
}}i`��~*�E�<o���.�G��ȑ�<��J�:�݉��̸�me�#�V�ns��,r�<wK���<��CR��6c���p~�3�=�����5 %�C�Wx����R)��(r�4�R��r��C�;�����^\u��!���v���G�ˈ>ݲ��������5��Im��l5Ď������;%5�,���F�}��mb��|TO%<.+Y������d�X�����.7�uضd@i�w�9U�Q k�R���d�D��w.�\o���(�9��D�����R�[�s����1e��LH�,��2 ��Z �܊�q�Y��tn��J��K[�ؒ%m�w �}��f]$������0���*���9p^T�PR,��an��|�c���[�wJ��8H��
��˒�,��(R�(D����/yB�{�_]�MnO��:v��F��̾ځ��2jJ6lp��C�2+1X���k'ݕ��o^��#4�ݯJ���
�#�v��? ���-��ѹ_��Ob���z�ЏXXcFM�3#O0�*��*>lw80ݿ��h�I�}�r�U0�� .����~;@6ѹ��)��am�
�W��Or��s���d�5���Z ��ǻ'2�=&�eS�Ec�	- ��;T�4��T����N�B�_�6�K#�ڻɁ�}'�B���؈2��KNj��<�p%ҙ��0 ���7��	������/�SS���"���k		�R��¹�_q��߀�I�ꮥ���w^�oV�ȩ�c�'i�fd�<V��9w��KHd�i�D��Ff�6�@����Ky�����A��Jg���_�i:
��؉(�d�2��4D��U�_�wx~�&���1~$J$�O8_Uj��SA��ge�`g���'I��r&p�cZ����&�HԢO��jF#����ڣf���O�^�,3�q��O�?���
/)��?��������LWE��҈�ӝ{'�	U#u!}F�y���P�=�J��0������x�~x�Q,�*hB��DW��1�a�{m�bK ���;���H��n��6�����&��<G��9�c��"ڤ��#̑�Tkt~�`��:$Nh�K{&͍5��">AŻ'�xTpH8��A\}7��TVL�$���0�t;��K^��M�Y# j��(�9H@��ʉ���r�#t����|�D�`��ttǿ�f�OE���J�?l1x���^��\h���s��~����HX�*��,W��xb/UB���J\r��ש�W��qĔ�O�̉��mb�kgy��iw����^g�|�,��H������9��E��9�8y���g�G�3���������3��-�E��Q����K���=P������Q��&7~�;��D7ը��O;[�ظx8bP㢷a���>\�?�c�c�y��tt��5��g!����$��\Гdf�Gr��?���vJ[b�V��� 6ޤjM�4}<�}
���0��¬QU�_�1��K�����e�!o�P@ն��f�4��K�EA��hS�Ǉ��+����{UΈݤ���Hr?l��m�1�mf4.ft���n�*L��?H���k$A��j���l�"(�	[s�C1A�.0�>�q���,�T��ٵ�8���kQܬ���44u�)�1�\h�P�0����eU�%&ƴ��l��:�X�S��_6vݡ�;&�ɰ�@�,��-d>�7�Ɛ�v:�e�?K������`{%����n��O��z�є|}1զ�a��Q�&2�Bȝ��<&�gv�g*Y���]�`��0��U�����3/p���}�a��l�(�����ذ�������} ������| N�NXұ����9�t�m��W�,4��`G?�T*�'����a&�Vx:Q��Y[�.F��nl@����NI[�L쌨9�8�* �xC��N����]縵;h#+C[��!W��2�@�s���i��������"R�o@b*�P����0�z��I�kde�&WkR�k���:������Sx7�3���MX;F<��/��+87�O�㎌���=���w7pG2ZT&�����-�`�Yf��M��	�7(��bu�Q�'���u�+=cݜfƞ[��q?A���M��O��+�j�M'�t���{��m�)�X*P����i���[�O��#���\�,G6rf&��T�wXG�~�p2W�[D�q�b��+��	O�h(�����e�9�ç�$�d ��Ե�U��<緎:�'{=W�W��M�J�O*���K[�i ����I�r��*�8�O
�L�)����Uy�Ɲy���NPh�
X��+��s���.>��V����BD5�Q�����+���\\��N��YYh�=�ZT�2vCO�'�P6��xx��gD8+�r���EA�y	���9z�U�z=U��O��i�{�U^&�i����B��{�.��ϻ������<�N�_h���0p��%�1O���I�o����6�m@i>�בr|[�3+>�W�4a��w����m�T��E�(>!��/�Xs#��� YŬF����*ȅ;�!	+�'Qt��*CS&���:������׷
�T�DW=�tilȘ��ND�XC^�T�a�ԝ�ю��,P�eR��������d�-t�Ŋ�Kn���4B_I2:�@�L�B�n"�o��G��h�Ɯ+0��D�=���J���M���`��Ddf6b��!�������4�\�����m�RK�4������Ӊ�@w�-`�O��l|ٌa`%�X�OXO<�HA(�<ƉV�Mv���*)���uLҊ|cW�s�+�I*�̬8��ϫmF#ш
�1�˙h����H��<,''�v��o��ּ��^�~�^�%"a.''q%��/�CzU�ʅ�: ��/�Q���4�&�t63㇆d�/���2&�Z�Ї:@��D}��ݱ*nH�V��DKf�O�����#��R��dHB�̻�e�����o�I�4�e/���6q�M�������$�uuZ5���-A ������  \��E����wz�lY3!�������aػ9��n��E��C ����"/�O�5��@5DZ��E�&|c���m	��o�[%�p����9?��R��r�hMA_���fC�~p`��#F���:�6�b�{Z�ڪf-0>#��l�E����G�"T]��ďP��7��_���a"4}�O���pL6F5�@mc�n:1�[��-�5�,ɽ1\� ���s;�N�Y�$/�?�D�[�Bk͹��s4$P_.(-�ץ�o�Z�{\�`!5�˝;5�!��PRlXI@�B�����������B��k��$�� 8����M9�3��pvp	6�����WU2,eПB�(C��>`դ�`��dU���əFza��g�I!hC!!����+B�|�6�qo�)�Q�k⽥��� ��o8(KN��o0I>@�x�����(�-�8} %}I�7����2Ԃ��V��K�Am��[��)����dC���M[�0��7��ݫ��AnA�5Ĝx1�`M25_�zD��g�X�~:����6K -����E|�@���]�E��z��;aAc��F��E�3{���7b���������,���Xl�iB�O�� ��0�1q�Α�zpPZH놉���Ȗ��ʿ�S�/�.H��a}����Hb 7�
�=��^/ ��h��l~zui0�vFV��d}FCٗ���D��˩�07�̫mԬ#�n��f�L^$�#cRlQ�����_%����D�����N��'�Y���M�|]Fق�K���;��1t��o޾�`0�CO
�$�ꉳ�HY�O�Q��>qiq���ż��]TH mM	p�K��Ic4Z���W�����噺y�������7E���)r�>ބ�j=���Ld}�e����~����ek�7�����Is�b7�L>�)����s��Ba�	v�gl���ר��P|C����v%θx�F6�n�-/�:W��V��O9�r)�	�1Q��L��q/�`�������0��fP}��A�(�1���j��l~������ޖӧ	��ō�R�hWk?�#6�Ig���z�ķ�	�i�w�x����Y3������Y�n0a��9)/�2�^���	�}��d��xW��'(wB]���^��R.%�.�x�����0e��x��V��B�q��������_L���&V� ��H"}&�'��{'ްM�&G��w
�
�k��XS��p��`�4~[̉*�\-:L�0=��+p���ELoxZh �m��"���*N��������22HY��VsB&<	���źgO�oyQ�8K4�u�b'��9�޳�<��o�O���t�0_�b6�((¹�"��?�$��˱�������xI �+������y�rU�|1�����4�%@��r!N�8^5Ng�v��^�eu�ƒS��5�v�Z�0�)goa�"W�w~߳i�R_��$�z|f��8�2���p#��7B0]d��L�Nu�I�?����2ˏp�dіA	�i!|�۝���#�n��y�3�y(��`}�-�# N���nW^�C�Y�k]�
���۝��߯��h|~e��hh������jS�wzM��ʶ�;ɸ���"Z�~���	=7��Ղ� x�D���8�m<��>7����S&�r���T?9��]S��~bz��|�r]�K���R'�E��@!Q���!� �Ӵ(� (gU�.�.Uم!f��G�=#��5�\�\�f��߷�@"��V6f�@�pP������� 5�3j����g���l����~��R~�F���b�h�������!,���/�Ƣ����6D�A��sCN�uKHJ�[z��a����\��HKy	Rֿ�7�6���%Q��b�33�x���m[� �69���_������Û���3�0�G�����X�k�L��P�<\v%؊pvZ\�-�����+^T
�4b[���Ƃ"���C�˕+��g,�'��|� ZTy�����Ы�1�@���o�p��aR�!H��y�a��{tf�u���15l�*
`9����M�w�w�����*������pos��@���F/_Q�3���X��^x)%d�-�-̴��N���gm�Zf� �ϊX��y%!i��u=�=E��/�Y�dЮ�Ү�.�>�L�՘0�RڀE 
]�1RrP^���[��̟)h-���%c��RX�zI7�ni���� 5�o�JEɥ�3��P,�B�Wr}�A��t�������d�j<�@����j'�A�DZ7�ms|�Q��n�d[���k��K��n�_�9T���t&���iķou�c�<��p�^�C	߫�Y�}
�����%��d�n�����NA�?p�t��t�������|M�E��>��w[3avJdj4x�L-1ڳ�5#
ʷ��éo�Χ>,>W�0J�*��c��(��B��k�����Z�}Ĳ7\}��4�E�
�y�ఄ��� �6�Qq���_���_�y��.����-��0]�ߞ,�/x�-�/y�1�\�D7:7��ҡ��i�jšx?�G�Y����^��i��%��������{�Tdx�Pc�,s^j�a����+p/�!'�J*�'F��aSm�M��jjN@��ꉣ��ޯ��������ݭ%�|�n�gW��<�@ �"�A�����x�OS����ġ!`�N8��i�ř+��������&��*"'O=˶�]�=���*�����5|Ħ���p�N_��Uo����*q���T��i�Үy�O'D�O�\E�׫̻�`%j�1��Ǜ�ܠDp�	��!�-��f�%9�uw�R�Ʀ+.KÑ�4�NM,
�c��,�	[��BCC���5��
XQ)n���[p��V�nWXl�P�t��ۓS֌��k��.\�@s�r�J�<��خU���(�G)ʵ�DoQzz ��J5	�.�+���������� GYc�{GBE"�XM���(�Hw��<$G���t�&�/	UY�ձf����p�����b
�OKkݶ���Fډ,�g�+]�ʺ��ҩ�������8ՐH.�T�/n7ukf����xE���*��(��qx �V0~P�����U`N�!��z��m+aD�#I��Q�?�p��@`�gI��`���Ap�EN`e����!8�W����#�η~�n�4Ou�Hj
 Gb��s5�d����Kd0���hG�,^k@a����f�G%T6im'P`��n���|{�Vf��g)�v�I��{�`SvO��P���o���x�S�.��o�����KY�k��M�>/6�'
�V��q�6�0���!�;��%����2�>���/vΐ	����@�e
�.�ӹ��f[!W����hޙϠT\�#�����D�k���D�)2\��`QY�����2\;�3�1 2ƹ�ݺ!��0�2�<��X{�e����K]��Ӕߺ�w 4S#o�[�fV����@�d(�+�:Np<ګ��Iҕ&�>GU�A�
S�/Q;��³x���#<S��4h��ʅ�A��������y3�mz5>��I��?{��/�@����H1�`-$&��m�؈��\�QK����-�ｅ���������]��*)�5���I�r�|''`�y����K��Ut���P�)�������9��&P��S�SOT0 ]9l���b���Ik�K��g��a|���ۏ�Ip�1_8���'����G�)'s��ĕv bz`�`Z�ġy������)* �h�t�Yh��� [�1�gݽ�;�j�s	�30��I�� ��fS���G]�x�/��<M��Զ��6v �[�K
�7I���{��'��	��'�����y� *�)�!PxC��p���cN��~��+��6G���<���[��$	��B`&�Z3�	���eD5螔eKhB�:��HT���Q�ٝ��5^�L4��yOM[��.�̦E�iu[���n���/����'%~(�*��c���:�n���~
P�?wn�Fm1�l�̗��\ 	���H�{�JX��A�28x�x�La��4X�im�Js+ʯ�}�)�4e�ܐU^�`?���jzx�t
X�&�ݰ,7�G��O\�Hߣ�)��-	o����Q��^��}�Cސn-ԥ8�hjWԳ�~:l�?�� ?�Q邬t?�2p+�����]B[�r[��ہ�6�ג���b\��ϵ#��2�~�r��ٗ�h����CM�i(I�u�̳1|�A��7rӌӉ�1���x��H��� .��.!<��SG{�V���}�t��{���`�D�;WlwA��𻽶N��o0 �Ɇ�3u:Z�h�z�.x[b�\g���@�[�|/鴌�E��P8��B$v�"���'�Q� �WG�U8��l5�ٷPs)F��gv؁x��}�Y<���������9[�#��\���`���^�]��`,�,�������]nih+�}e�S|~��m���5f��D� ��M*�}^E�Չ�ڨ���5�U�8~E:�Pf7��1��ƞ0�sA�5KW^?���[{�9�ӭ$�Nڧ0�Z?�&/�5��69�n���<F���a�i�j���XL���9��a��I��*"nxvn�z�z�-0[��dC�<!�O���kMVf�����H�!��s�M�f�Ķn��r���r��+��pƝ��"�D��V��_vu�W�F��ҲR���}�/{m� 6��Q�<��e gl��*�>�rx�� J�oww�¼�KT��|PM�v��)i�"�i#!v�����ݒ���|WtPs	��r������s�JM�
�y\BJd�̧������ �z:&�sF���z�\ ͧT��KN�{�qH:�B+aޮD=�ƈ�0=��������2^���	��_�Ķ&&����?�[�x���f�?�*�q�-4"�����u��ڳ�[s2V��aܭ��95�j[�ts���R��@גJ�a��XVք�f�u#~DQ2!	*�ܜڔ`s"gl�E�"��m&����C<Drz$z��sf]r!�s7��u�����~�C��V(�46������auw�b����ro�����Ke�¾脗R;����I�h�^��2���L���D�2�f��݀3�p�"�J[`t~E�F��
3��V���1eY:p��'l8�@�y��Ю��%I;�ε��ZÑ�FgW8���N%i�
�\�{�~W����j�|��?�~SP���b>\�w���Im�Q�kxC��(�,��a�e?<3��C���G�n?W0�<�cf��9{��Z�#�؆����P���ӈ�2]�˾��UL8��s�f',A���sAG�!�ȢF��CN�:��Ѥ;�����B��o����fG�N:%p]4�n��P�?)(��'sj��'�������=O^g�c@�ʲޱx~��@-�zEV2�� NE�5�%6C=*���q���_��2���W�F>lv-�яn�{�l<P�"�\�Eu��,Qf�7]�6w��E?Q�u�M�����'��=�{�K�TO�%gk�,�~��Htxf؁CX�Ð(����Ks U�cR(،u��r���P��S���H�����X�5m��Lt��!dڊ;�h��=��&xK3V
�����L{vLM޾�c��II�8ɬ?�D����v�,�B-�L��S��N�U�ǐaqJ�f�o������R�=?���<�3����|
s�~�0\�;�Sn/r{@n ��@���]ze.r�5��-P3q�|��ߣ�y%�l�j�D'xÞ�U��a�x��K��-I�~�4�h���Q�D~��9�	
��^6�<�R�|7��S#F�\��^��n�M�t&��>�E&�����؆?��,9zk��V븙'�{�k�����<;��HX�;Zk�v���<#96uFh����K�x� A�@yT�Z�e+$�������M�C�6r�g"�'!EX�#�U ���?�NV;
FP�ӤG��<w��և�"�\�8LȲ�b�K��Byr���=�/�,����Hc����[�1TH���<8^
E�r��`��a��S��XV���1*�}>�G�#D��o1���?��ϴ4.Ue\�)�1��rp�tVl���ʑ��8�������wX�2��怽ד8{J9�
c�O�aq�[l���b�y�[Y�œۓn	�@�i=,�j&j��d�Ub���^k�37��S���S	�S~�ۧX��6�`#���<h�҃$�1c�	��_�L\/djI��؅e����c��w-��u8�RB��bY���5�7��N���F��\�h

?_��n�&]d��=�~�}�ȳ��:Q{H���+���m�f1�3Ƈ:0��m����(��\sC�)��W���EH�=��dTu�7�%�z%���X���=�=�  �r^��?CKP��-�=�~�N����/EλCz���[��t��ݝ�/#�'DH�&n���*�h�c��K��0qM9�?��x'����49l����U����ԟ�����\0��}z��!���y�а�j�������I�^@|��5�����Gfq�6_��b��H�,�����k".��q-�AՌi)��YP���j��yn�gm�5��xeV4�m���	;��x���{���Q��b���_�x]�