��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!��ߌn��-��,cF�W���oS�\7b��&7����p��N�u�25��D�l�W�=%�1�Q�jzk��Ŷ_��s��Ȓ��{���������
yKR��P�*��*�8-�A�)�ӪRG� �j~����:Gd.�TB��C�m���`�ʰ�l\��/-��W&�R��ѯ�OP2�>�Ƥ���]9�r\�~�-�7y��;7�����k������,��$B�0jU�m����+���x��
��\�7+^W'�o&��Wd�YK1��/k
Z�@,r�~��-���<j��hVhp��p�5�,+J�m�ɶ �e.�t4����������d���q�v=>rS���Qˬ�,D����*�8�fI���ȭ�VFj���\N?�Ŷ:j���צ^��8�ʏ]�����u���]! �J�$b�.&)Tg>��D��h,��e�T�{_�b1�_�ډ��5�Uf�nM���'�u2�$�����{�E�n�Xz����L��
>��� � ���	
K�υq��d������n������ˠK&vZ�Ɋ���5Wc�+�q�㘃K_B5�Ԗ�������3�ix�6�
�+K6d��lF�؉�4/v@�����Z~�K5�� Nֲ?x1�'#����¸�{�W��T,��%c<I?�D)��v�+�f-����S�G%tez���F��C��3t��z׉#߆��3i/Ж�J�7�Ԕq(�=1�A�J��c���55^�N��𞎋#�[���;�N�t�Ñ��_k	��qIAǎ,0a�u_�̞��)M\�]�XxV�q}Q{-�3uf!D�ӊW��%�b�����Ǒ���c�f�����V����=�Tk�������k�9���Cڝ���:d�[ y���c�Gof::����tiŋ<��w=�j�Fٳ��ʞHe����q�fBy�����!�����J-����=[�ĸ�M*U��@�}�H�x&qLr�3<U˵7�QI8�*Y۽o���_�̞�)�B((������!���>����S���LT�R���z{�$�\z$���=Sæ�����o�G��=/��/��'HҰ��$�W�X_�yQ�ı���?MĢİ��E1_C�U�E��Rh���}7^
�w|�/�gt&R*�1����Ux�OVj2��h�O���!��>�3l-�K�T�S^�
�N@y���;j�Z(��×b�Hޫ�l�(����n$=^X�W��8�z��J,���(�d0�������_��.F�����Kc˥-��|,ɵ��&���)�XD�^�3{@���AX�Wv$�V��E��*��җ~�2*��,�BYxO��O�����~N���\6�J�h�VQ�t��cD��pbn]B��n ��0��>'�yV��� %����o���:��>��M5_2r<�S!��w�O�l�}��#��iR�7�wk�R�o4�U��A�����&;��V5N�� 1��\������`&%�~��0���=�X��y#�>��ZL#b���ϡ�YK�67N��:K��w���% ��������~BӜ�w���f�0bڈ�9���(J�@���� ���guƕ2��wrc*_����=���i��UA�K��A��l�u�m�g�V��Xd�����*����^W/��#Qi���Ψ�58\�k
��~q� �
��n�C��x�hy���o;��4�k4L-�C0bG;��E1K�0�A�����\̷�8f�7=yh����Ykt�U~O�Ԧ]xg-���s/,y�nX���;,4 6ߐ(��?�@�*�s:u� ���9Rĺ�/2���.������C��J%Hj�05ϕ0wԈ^0AI]'�d��[��ό�Fž�z�p#��(���]������;��Ͳ�@/�W/s�R��(d}�|���'`c8��)��Q����V��"���{�A~2�B_~�2ʹ�����I��a�U�M5�u6;^�{n�ˢ����۲*7��Y��c�[��(�HBj���	D�-ԓ=�ͤ������u��g�qaX6k�{�b-�.��x��	����碴B���J$�#���2��*�eȭI���xl֎��.y�"�3V���+\_��p��b��p]C�C�@#��}�2���WF.z�JD�����K���l�qI󎀛 ���W������OΓ_�2����Jo��l�Fޫ��#��{��jJA�zJV窊*�Ί�i~u�,�����I�y.V�s����Qϲ��	~R�pw�@�1�&�c��&å�����$w���nk!�{Vj�αX0�!�s	,��v͢$ɢ���f���:B��n�)h��{�Ā�G���O�v�I���j�������ծMЗ�*�һV������5��j�Nn1����
�6������7�`\�ڲ���9���Z�H�M��5a�H��,�Vo�E�n����$�t����%N��9�l�>�4�putG��S�MQ�u�sc���|�0[x�)���� ���Apn�0=b��Xf�$+�0��X9p��@�\�+E�m2�}i�ɼ�j���˝��
C��sZ�j���O������J3OD+��;ua��%X�@q �FO�����z��ʰ��]}j �;z��|^Z�ӕ1R�?P=��l	�PR���b������G	6A ��ZJ�e��,̝�D��-l������<�7��ݳ)���M�,�F��L2!���n�S# [�k�e-Zz�/R.p��A��n�۩�KyiV��{�����ÍtE��W7NDU�� #�pPV܈�̹7��f�P1c�C��.dr��i8�nd� 1�(�����n9�����d$����P'	�I���e�T(?X��e��U�[Byoe�s%�wQ��ʠ����?�{��*���
�Z�ʸS�t�w�c��#R�cѧ�s�Y�k<�*�/\d�s�� n�0���X�A���1��b��v�T@J�xb%q��X1�>=Lj����9:�48��O�����:�`�xl��#���(&��s�܍ďwp5��R���w�T05$Ց�U�10*<�]���
IJ���o�=�ȆW�lO���M�`#�)�����=gZ��=fZu��R	%^{�(�g���⭩h]]�>@b�k�|9�9{ތM�mη��݄%M�(�A�gom��e��ipr�6�� gh[,�kW|���e���#��e������A0�sU�ֿ��"��oF���wUp���Ŭ�>�4�B�{��qĂ�~3��m�/e �Yqt��Z��	�&�Y��x�c���w�ܱ��]	��֚���W��*nx�긦��UNѷb���^��Z���i�.�nR���`�����$I;}MP��a�e?x�ә �voExE3���:��Zo�jz����7��G��']ӡ����QO�L�){#�P�`�]�"m�WWj�� ���"��P�qܦ���m�m	b!m���0�9e�pD:�\S�C�s2!+�Ҵ&�ck���^kC'����mn#��I�ot���{������٨[?��)/��B�3��;�{we�JHl��\�P�6�.�+�Wǲ�YȾӧo�|�:YJi�	G��.�+/&Q��0(�fA��+Dw��� �򠡚^�2��vg�E�v8��p�k�h�w��wV�yq��F��UZ_8#��1���;�5��Q%ܴ��lV-yl�q{��g�Uj�q����C�����_�9���z�I�ʺj�Τ��cB�We�aa^�-Fo���蔐\�{��֓�
-Ջ<�i���0��=�9J�Dph�𹴄��ׁLQ8��ބ��7Gs
�Ћ��m�A]���nĕ�p���ʪ��6��=훘	��EM<-�M>A��נ�K��\�U�j~x��~�Q��K2Bh�םĎ�q�jp�����P+�t-ڕTt;�5�V�Lo`e��A����e^V��/Q3�����u/�9���rK��<A���L��p����$���{�r�us����x��b�[]�� l��?�϶,�\�-P\Xo�r�'���fYqn	
��c����*$N@��N�w$�	��m��n���:|�o.ٷ�c%ݶ��Zр޾��܍?��s�}�Ռ��'�	���1��5�����s���/Sӭޛ�o	G��%���}�N!e2k��a_י�$ʀ��Q�t�9 <Ǔ(k���f�[�ЬC�<	��AG`
6����ng�Q
�D/��Z̈́���˓%�����,����@��=+_g��Mt�@��xu�tW��M�&W9Q�Vbv�o#�7�;�QJ�Ծ}���8�ʚH�<ၺ�b�3���5�$1�����!m��\�@���xG���-z�������	K�բ��p
L8˚ַ1�`0�?N}���U��c�P}���	�����t��Y�ߟ#WK���Kzz�l{WBȷ���n�hp7��D���P�W�����Z¨ΰ�s�Db2"jo�4�\���r����>>@�u-/�]�c��Y]}�ɀFK��K��~��G�0��<�����X�sAwct ���Z�%T��Av�a�'p#��o��}�ó��}�@��"ܬQ�Q�����b�)�� e��YDqWE�7��!E|>Y��q̖��#�F~q�hḘHӅj�<�{�(L1��&17��|M���a��4hQm&{���_x,������i���s����Y1m�R�ksɣ+������پ7�������tT�Z'��A��E�r��O��+�f�Jp�(��fO�C0"�|�M�fF'�g��S��w����U��o���aSD�PT��MY߂��bQ�E����?�m�#�]���a0ܪL�Eջ�E��"Q"2�V������B����*�]�׮B ��5��ȷ����٧�/�Mf�����q��$�Uؒ�	HmK�Ti�]��B�������7a�������o���l�1AD�
%6��]ָ%O����u/�?��@N>�W���C���Vݟ��v�|�\1�M�]�-<9���x�M��;E-d?��խ��O��F����������s��u��5w�1r��m1�4����ը��E�I�\���o�Gr�D����$P��q`�b��<�X�䳵�ӽ���Z��F��j����(�O���lL���5���PL��L&�'��Rv7��u1���_��pR!�gԼpw�8�$v��K�X#�ˊs3�jec���g���_�@�8xop`�k�}{l���_��kÚ�Y�r�5���k,P$��L5�ȿ�?W[ƞF�$�"(>o��	��}Pl�>�2>^/��c��5�A0ZD��&e�ˣv�#	��S�ImP����1�����煊9ŸN��J[`�"1��#���PV>ڸ�&�!L���I��8�N����;'��.Z��(/����%���{i�P#�I�
�+�i�=�0@iw���I�,�k��2;]�;"\A��8�;���3�n�Ώ����KU�@仅1c��JX��X o�O�`Ia`��mhE�e�W�$�i�.�}���C�odm7�կW��e�4xU�EDOV�yHo���m6�''�&��#Аv���U6������ի�Ȭ�M~yW.Q��1?�}[�9fm�K����C�����d�;}�3F��t�I�+�c��c�܃qԓ����<�3"h��|��6!����g���}@��c��\��C�����+X�r���b�͜I�W) �(蟱)QF�s�ŏ�5,�k(#��QRJ��-�x�i].���0��WJ(��qvi%!���n� "ϧ.R�6���I������ƚ��9�V��ڥR��65H��G�^̩Lm�a�u�5��%�
E<Ru@ ho��@B��no.�坉ù�	��RHh;��q�ᰦ��L�i�$H����ʛ�"��>�Rn/�u��UAh�� ҝGߧ^]�%�V�ܪ���6:z��NRg�I�a��G��Ő���B�.!!����D�K"v����u�	M̠��N4)��dd�E�S+9���`-����j/P�R�y� t���7�ɕU_�m��^��3b�_ϓ����^a�/�UYJ�J��U�D���45�N�}%�晱������ <0���{�qfh^t�*.ԣt�8ݹ�b�h9����Z�Q#ق����YςO$2�	�tRo��¬V`u�2��M�S+۴ϒog�3<�����J��E�̴ڐ����p%>�'�f�l�κ��z�%���Uk_�DG�33�Y3���e)ep�����eЄ��*��RR�U�y&���UL�Ml�����؞���Zl�͛ъZ�m�{Ioj����e�e�[���:>��~�?�k�x���8&��#�g�;ؒ&s<a��+�o{�������<mW��{GO��_KǢΐ�B�H�X���{Ḅ������غ$?�r��N���L&���*1�Oy���Mr���R,X!h�@������Ȗ�^���ȹ��ņ�-*�c���#���̸cs��U\E��GGE\���Ѵ��1?�E=f����0��yW׉�L
�ͣ_9�B�Ke8暠,9;R�=� �2�z��[�G|��-�������`Z���=�&���V/C:�����XB	�όK�c���P�����+��'�Vc8=a{�L��y���j�D#�lIȏ�ڀ�����`�˅i�����+�1�n�Cu*4>��l����ĉ����-�BUP�ŬP���p��)���G@U�������"��UF�.?��q���������jQ��C\��x"W"�����;��D�;��;���|�Ķ�L�#?х��٫>�Nyj�x��Ә������_�ڹr�� �A�k���P2S~䋒��o�����i�:����?�Ç��̴LJ�
��Y�����:eψ�i���}j�x�r4b��3�`1�;2�-��%I�,����c�:Ch��h0p�j�}��>�GL6-�8�����v�S<���R�������Vh�s)�Aiw���0z�F~�^�x3�+�,��yz�UP�V�S�,�(V>"�ȜBd�B׀	/��Q��y��hّ���k���oȷ�L���>W��^�]�c2FZ�x~����=B���V3�X�ӆS;T�ڏ[�=��=%~M�@5U Z���7DU����3}3\*�p����~��2g�*5-�/]��g��\Re��*�#L�/Ui��T�Fu�фn�A�ѣTLh�rh��)v	���Vs�scЭ��o���7
�^�,=&�}���J�
-�w=V�H���݁b2�qR�����ѫ�U�k�Nx�{.�y����tm���::�<��^me��4��.��	��\F��� "��Oˈ۫Jzqp�gN�\��fG��;�\�䟟F��\T{��26��wCyb>(�:w[��9Sׁ#�wM����a�^y�ߡb�kk����z�mЃ�4#�V
d��o	Z(׿�e;PW�ueb��n ��Zh����E���>���Y0{��@�8�Xh7lOkϿ2���ְo$�S�2^Y6CB++8M�	l&�4��n�.�@�K���< Lxs��k�8<|��� 0��]ow��{#&n�y#4��,�K*��/�����nb�pן1*F?��5#FP��϶��l�D C��lz Pg�P��V�֔���X{7.S�����c�|�-�*��)�u���_�~�f�@؈I�TG6�.:���9�I;{ג�n�� Y۬��ùGۖ�7��B
`��7�8J��Y�p͝N�g��#��=q虎R��y(r;�r�ktR�5��]���?�Sޞ̈�q�:���<��w���g��5GW����i���u���j80UW��/���?�5f0LӪW���5G\2T�D5N��pA��?�w�v;���ϡ�%���V�e���5Ǽ�����F<��uC�؝�[ʪP3��א�X����@b1b���?�0�9��).d<!d�����X�F��N}�����Q�_-S<�5@��;(;�"�[M�%�a"J�K��МՐ`)+/HZ)5^d(V�T5�5������A�̔�R�y"�}����P/�S����=C�?�Cb�P�-�֮�}T �B%$�ISHS�:i;�.��^���?$�	�����|ϰu<�Yq�=��2E%�����:X$�ښ$@Z��`��n2�E���_V� ������ؽyѮ��Ě��v����*L5�YI��/ 		�G����Ǖ�F$�4�aM8#n�%%�����dB09 ��Y���֣�=��[�O����%����yO��i|�->�cd<�h��:��u�l�Ξ� y����9�H��?N�� ����۞�F�p����{C��͊�i��s{fD~� �qvݝ����񿵻E��6��n�W���2	�M��nh��&(��-���D����R<��S�>������~�͹(�f)Q�n Z�8vݼ���Hogu���ú�R��.��Yf�O���������n�T���z���=m���_�#����V6��*�攰�l-���h��gTx@��8�u�4D�н\��
4����T��
�"�c�us�P_(w� _Y��D���>�&WU}a���J&����X_	��j)���^Ѱ�/=����j�g�$�2?j��
��K�����̾Ѡb�V`rk#"p��ML��O2n���n$=H���W}͞�źƚb1�RA��ap`�1|҈XI޹�C���V���S��وjN�]�yO/�:���0{?��Ae����?�@Q��xzFA(���Ѯ{�i���lC�q�-�*���r�nÃZ�z*�)\;\#Z�Qu8��A� }��&'��߾T���l���ϸtT�s���+���~�a�H����F���~k��W�/�RΥ�q܌�U��+�٧�R�4�aQ�יA���\�j�Ly|�RI�uo��El�6�°i�9��S`��Ky>H?TMy��UIyA�f{�=t�&��#BZ=�ٮl������`�R�{d�s�Y7N��d��_:�g@)$�8�t�ˇ�	6�K�Ձ��=�Θ��v���s~tVO@��#+�f��~2��#j��m�'���\�K8*��k���r�gZ���Q��C��ZMNy�[G�k��G6F��ܽ��>�[���]Bõ�t:��f�����o��ia�6�v��\[�n��0��1�?��Y����%チ��-g�C��=�w�l�P6g}�ˮ��nw'g�B���Aب�������ٜ1ڵy,��,���򀴵,�����N����+t�fIfd�wK�'��=ʖG���������j%C�<�/�䲆����S3��X)�����S�W��__�o�~%�L��2�Q��]��a���ʱ)��hHu'0�٘��Pݡ�ց]P�藁����k�cYԻz\Dؚe�_}֓
�-_�{2����\�6J�SH̚��;��<�f�R�B}>�-?X��-B;�E�0`�A�O���F��Z��:����kӒ�K��|�\^�T��5�t=]JDhp#�;��s�r5���\�%a�ſ������l����~]��y����*������lxA$�ϥ'�VЫUA��(_����i/,j� ��Nd�4�bP!q<qU����7_��-/�QUJ�gY�e&��,!�mj��%��^e0s��F��O���C��ֲ>;N=3�K��� �=�������_y:Ar𑻍�T���X���pƉ11���&a��ZH��f^`E�i��n T�`s�p�2}�@�ɇ��,L���v�q��	F����� I�\+/��-��+u��-�d��~�yl�f���p0+.��w��.��'&� o�)t�J������59��G�^Hӗ��W5��^&����O����-��7e�79_ $yck-<��=�2��Ymw�0�	�f6E��KwE0�!Ȭ7c�.����;<q�����J�����/]�U����M(@����M��
��UޑA�?#�f���sX�l=���9qZ��(�Ә_�5Je���Db���#����z��"��1ï�
�1��׭�j��%��L*��ffÄv��~�2��	N��j�x>�ט5~f\�� ���<؎d.]o�p�{����^(��BفW���B��6Jj@�]���*�(��`dk9ED�|��q���jI�\��b6y�}Hk��J�r�3,���RV���܃�wir��:�@U
��;���<��Y�*Fi�zzP�Z<��Yx�烅6�E�F)H�
~@�`{Ƶ�/ڷ���M��+Y�PU	%|���,��;[��a�c��Z����Y}�j�w^�:��?⾜��#�|:��������eg��^�;ɥ6hz}��c\�2�\��xud����_�'؜=������n��6��1�O%Q���ݬ��A��]G���NL�)(�����|�}&�@�9u����_�hO�aK��]n�><y)�y����3Y:�(z[�?J'RTf�Z)�V���y��l�^�?���.!����e�lk-mǒ��(���|�vJ��T���YX�S蔨�������2�/9s���J�ޏ��pֵ(϶y+���YNZt��1�������H�:�*)&#@���</k�e(X>7��n?5��p�z�Ĺk�j�i��Q<g�OYc��E�	�A�
�e�K��_��7K!��Y��q��V���� j,���6_W��3�O�%s�-�����j��޿g�s�V��t�a��t��Z���[��~0-�I�����G�>I��h���U��n��֢9I_�=	w�/���@ K���~��
cst�S�IŻZB!��G'LC��%��5����0h~�ǇEJ�"�<�MK���؇�Y��Fh� ��.� ��1�(�C���XUq(��\%d�Τr����b>珞�ܽ9� dY9���~��*Z=�������Q�gպ�Q�TaY�X �|�0g�ը����H����<�g##lʤU�b+�H���$%]+?c�V��)1b����mK@���z�u�=yJ�9���B)�Ǖ��e�3pi�^�����Ֆ%��̭D�!ӫ{Zx N&��+�l������t���=~�*��N�)��X\m�o��a˯o�,�����9w�Ze��
$D���+҇t)��5`���*Kh��X��`��7�C�ń1�?f��&�Bf�@�0r�L#Խ�M<_��Wb��4jO�!x_�Ɖ -oLe�q����IM������:���?c:S���@V� �[�Ǎm�s*���`�{�.�0X7��H1�NR� ���8�Pbe�q�ӥ�{u9�иy�U�}v�*T�5�2����t�섆�W�O�N�Ԝ��:��P�~����H_׏R�L�v���"��o���1�
�K ��cRV3��t�ݪĳ},dH�-ʭz�T�t:���xL�J��ѰG]&?8:����Tꋲ���.�+�{2���wG��|er�ׅ{{~���{y,C��
���F�"W��`�~�NVf@��T��	��z�C�`�m�X�w^O���R�
"�a��V|$�d�߇�d�÷��0}�A�xF@Jܾ�~�I!�%Tg}X۱�i!}e}���\��C�X���R��0ß*OWf�d2_����z�����F����v���5�z�����ЁɆNi�3�!���ρ���bژ�A/'���g�^�`;�'�Kj|L�����﵊0X��d-�'+��,C��6�6^�"Խ�����c�*=8!�[���hܡ<���|O��2�	Ġ0t��>�� �(#s�¤{Ë��I@s����&��[��	|���/�BH}����B�䁈��GR�kc~ƌ���Y�4b�}�ʫ�T�8��㟃��£���?�.[2�K�-��߉Z |�����!>�x����L[�sc�!3�E(���msu�~Ǟ���1E�5���`�V��X��[��4�Vl9G>$�����sW	����\��m�Aa�U��5���8m�9=L����p1�㐎V�Py�#I�";_k��7^��y�S^������8��$�[x���6<�l��d���=�x���~nN���ߴ3E�`�kZ�Yzg�H�G��Y �,�4���,�<ס��cݔꣷg�C��`��D���W�B�P��7B��4�ϺiJ�drH�S�c�g�XP(�G�UQ
�ܭF���+�k�s�I���AsZ3�%��o�>�n�V�s:��`���
�_dq�q���qgz�ގ%j�޼�Ʒ9w�.��k�=��pf�ZC��%��K��Ym"���k�^�[X4^���*`��y��z�=E�)���}��L8'!�ɮ!7W�	���.[��|����l�-��n�%g�1֥����o2��:[PZk�.���|d�4��Q�P՘K-��RR
* S�����z~%;#�-�0�|�
�B��
4�j����C�o���#�de�L�T%�̻9E�1�v}����D�l�
��Gn��!�R0�`.�r+VĉD��h_F�(�����a,�=-sX��>=��	[��K)�2�=5<	���{Q�jm��Z����f���5B@�TXtDk:�{N�1BhCP�Q�Q���ٚ�����&㲉�Εg��.a�00A�:�#��͝����^?�#��0��yCLb��M�>�>�@(k�bwJ��iq�j!Ώ������%4�[=�X(���}�}����f_I)�[�fR՚E�vZ�&��'����*��\	�,�8�7@jO�M����ƀ��U�E����4�D���?j�v��w?������R����Ќ��U��t����*���Tǐ��q)�K�vոw�!z���'�?��w�_>�zzonA>9��[�b]|_Ai�1�|�0]/���m,M����2$�s˕b�n6K������5h���%��Ka�@C@T\�cV������8m�`��S�����E�T�86� �u����lax�C��3��zZ��ɩ��T'�r�vs�_ �� ��L�����g��[�yc��0i��V\'��m�D�4`��Q<`	B7�ª+��#�[�����-�����	Qի<���@ÚP��}��9ЩO*��~�"I8�x\Y��d��\�w����b����=��E�r%�_���Z,o[��ֻ�Xj�'��zz�$�\̈́��u�3h@(��h���_[�ȅ}6Iٯ�lQ�%[�=���8�� �䆃�)"h��l�&f6��V���ƩG��N`��K������I�E�������"����ݴ��Y�{��U2PPE��)���� �Q�~���R����f��MP��E��� cA=�ӽ6k��b�Z�$�Wt�Ŧ�������i�fw����	�<.et�`>�w�Ep��X������O��D�!�T1 �Č�~����T���M��z�9D�&'���6�hN�m�p�=ʨN�����]�u�Ox��5c`���	� 0P$�@���he���ceLK�������3�9{P)�mP�Tޘɤ|�����j���sC��*+ϸ/�OrCf�+ [.��."�����
�֪]x�g�uн)��-�)Bp>�q���X1��Õ���Ϟ�C�n�c[�X/�z2��tBK��H���tU��D$�9և!�5cl��sa�ac�E�9c2�s�g߯�=��V��d�A���R���}�2�O�Rnx @ק����{5s.-8]��^A-�f�搹5�c����ɢPxn�$�t�@��
T=�A~s��tSxhcP�yrs��?$��ro�(��kB?
x	�����v2�n�!�z	��)��}|��tD�ޏ�x��ܥM>j1y`����^,���Έ���L�t?�I�<rO�p��)���2W1
��d��|���^o�l���c�ZE��+����{�P'��U��D*��rth&|_ 1�ۮ>%�}ƭ�;�/v^z�����wR����\�t�G�}j�Ij1Z��p�:H<�R!jF8 ���:>I���F������o�]]��=k����ϻe0���Ⴘ�L�'�8#$��Gw/��Y�*���%)D���.�v��uc�u&�D�eOK��|�X�HN�%���_� ��K)1�J�3�����e�Nڣ�IP(�;h�}��p%?(�x-jy�R���TL�؜�Y�9V��M���0H���w�*�f��gz[%��h.�����3X@#���(��ȕ�'� Ғ8�:�5�ΣQ;J��luvs64r֒{ػ��{��q06ߐv����8��z��S���c�qh��E� ��*�����`µY_e�������\�P��'��>��k��'�N@؏L�Ľ&V�;�q&!i���.@�<���Jt��}j a��pW��L��V�Q���pd��τ��d��O��٢�~��c�"C��Tf[�����,Eqc~�r��sef�%�T5����lߒ�۬���U욡=Js��9�#A�B���r>�L�bێx��+�y����ܲix&J&��� ��7�P��`ĮG���4�2�����l�r��$��S���?�ؽt�M��+�ڴ���of%3!�!�%�8�Эt,���z��4�7c,�y�%���<��H���ϱ;�ힶ%>����׷�N~�ӢK�Vf���L�.T���������#b��������eZ{���w�d%�뚇w�.K��6�V,�)�O�S�����,��M�K·ׅ���>2|��"����#��P	��2��اKl3k�61�^Fg���gJV��1`
R��5,�'L�E�zk�g�9۸��r�_G`�fFxa{�N��y�
zƤ��ګ�"?m�n�t�!���^q���ݏ_cZw��b�A�j�H��Z�Y���5��r��.8A��ɮk0B���F<�����j����ցfz�0���a�$���Z`�zq�Ef�2�t{�*
�l~̓����i�5߸5�E!%y��4l/��X���z2Ə�L=����z5x$���-��a)�_-��h����&ǘ��"�����2h%i���F��)	4�R���MQo]��3�q�L���H���[���Jt'w��D�F��)7%u�@�g�{�!�1����8���'�̥ ��6��DW�jDG�غ�Y�v�E����Q"��G)�q�4l�ϯ���dRv&�o�
���]�n���csV�ڮ+-�g�E�X��(��Ҳ�m����-��/{3�Z���6+�Aq,�@��,���o}��e(\�y��{���m!X��A��B�7��=p������9����Kw�
J�]7b��nK��[GZ!"��m��A��'0�(3�n=����S�y��z<����q$-t'ҷ��~�����t1w]"�ւ�qb@�1M��]��QӉ/i}+���+�޷��&$ǰ�[��_�T���q�A��$�5��BKW��~�����G���3p룥�l=�ػ�B(��Uf�5�M���ӟH����#��Ap���˵��V7)u�jՔ�WV~�=��l��r]����x��<�	��ٔ/nOv�Q���͞�_�,�V@/x��o��zn�_9����[ 4bُ��mxx��i5uȪ�"���;
��4���Ň�c�&�-��`e�܅{�E���z�F������'��C�����:Q~�}^�7x��5}Pq��ֶg�Sd�Q\�B1C3*�lg	����ƑJ��V��B<+K�	1���Ǻ�?��N�,� �N�Q!��QS�4��S� {�琪��b��<��v!�h��bVJ�Yz�>��p�V�4ղ�ߙ��n�+C.Z]|̧Խ9�� �0ڈ�L e��l�R��h.��c�1�G�.�%x�s+�-�N��_����G΍1��^��=�? ���8l˰`*:��J-�^[��j�Is{eG��^�W5)4z%��S��վ�;�"�/aP�G8s��p�=63�k�h,����ԭ��3*��g6�|��y�%
��Ѧ�'Сu�ī$b��K�MԤ4ܷa�� �lh�	���a����-&�i�ΝR���⷇yU� ��d� h�b,��ʙ%{ۥB�I�AZ̾`����S�_�OH�c1_��0j�r�#l�	��y)�% �k�d�������	RT~R6З�}����'r�j��`"�X^^q�җS?��$A���:������E�l]?T�!A�ٲ�"�OP�lI��q,������Tk9,Q
"ζ�
F��N&�����/�i��N&� Ynj!�]���3K�y��S��)j�x+.̶ϊT}��x,���F2~�R�� ���m
�{��5���o8�Pf�UDB�*"m���L�zj�9�-8��.��W?�4F�ɴ�X[=z�9�w_Y߀6�<g;�{L�3�:��ס�R2N�CF�q�o�D����������Ha.1��6�����큫�����dȄ�fQ�-�FMU��a��EK|�p|A�D��y$�G�3Nt޳�RT�w�ɉ~�9	%�VPqءG|�R�54���Gp�G���Ӿ�6TP��<������;ͲwY`}A��/p;�*8�̟Mߐ��
��Q�hJ�X�`��q�����O�M�q=�\La��v��l��ҴSe[O%�=�W�`�Pw:��u��[aF6�`�X�~�=��%1ŷ����8��4C��$���J ~��"��Zd���X"м�;<fqe('�D�àvc�F`L��ILBm jRj_z$�29e|	��@�n���jX����"���yU:3c����x��c�)r������{�{V��#�;���� ANUK��i���87�x{��0�����H��l��a�c��TL��p���4���1���E�S��3A@=��Z?����Aڸ�
�h4U�?��:i��_�:+ֶi<��_X���vZ��N�"\�|�b�N�`p������c�ZsЦ\�� 0&�Ϗ��V�s�.l�w�a�ɍrxU�Ľg\�6�{o*��R(��#QV=t;_�ף�AJ$��~F�n{o��Ѝ�UVQ�N��%|S��
[��%oU��5��9R�XPG�� �ZT3l�K�Cy�&֋�&�C`�T��H���T��Ì���܃ʩ���mP�M7DU��P����gm��VƷ�
���N�.z����-��LY����L�����Fb��I�N�GU�nZ�'�4���"�ׂ6����	��Rz8:�J��[�X�Ѹ�b���,ãA����N/���dP���G�p�� :;^��7t""j~�A��Ϯ��у�2�U��t9)j)�M즚x���� ��k*'�̷��}��N���{	�-,֙3_�즷yS�������&���~=�d8m��D��݅���q�]��P�r~7>n�M$U���M��+�"F�}���[�n������g*I���P�X���J��G8_PZ�_L�������ȎB��_T��f���t�w����i��� �u��`��aj�̂;��}�j{��a��H�n�΅�	��>1Ix��D��}�E��ɴh��[��Ʋ�3�kY����ǕÇ�~����Ųu���f�5�ն!��w���F�u�9OblϔN�:|�b���D#R h�x�T}I�0g�d������\E��ǭX�Y�t�j���̤ʥF>���l�����N*x(-r���a&�o�|�X�`Ty}L�R~�P*�yS������h��]���/Z��Z�)���7N5�� L��2[������ˑ�����S ��8c���v0/!_���l�nȈ�N����>��G��&U�_�&�_��vZe�3���NՙT'7gٕ������HPwZ��;_���:S�Z5��,1յg�+�
Q�mdw ���H�yXa��P�g���F�/�����j���mX��>@���j���Nj/Ǵ=��Ő�OC?u"�_
Ǟ��
�6>+�8�L�[!4��l$n&m{(pN��{ac��W�ۗ7:�h��� �m��A�i�<3O*Z^��9�2�5��^[