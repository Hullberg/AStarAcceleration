��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���q�����W�E�9 Vοօ�̷�S�;(B�����",�U�s����6���i	t̂9։l�W%���Hl�1�iS�S��
��.]�h�9�?�s�_�~��� ���"D���ԛ���,w�K�te/��\�W)�m����Uq.#���,�#�����E=	]xBP��C�q[�������f'�H�f����3Ar�mӪ�������Zj�|���;�w��H�;/��dey�����M�:�'G e�Z۝ᕶ���ƞz;��������(�#?�a#!aI�X�&��G`�G)l���U����ս��Վ�8���c÷һ����PD
��΍e�*�[������o,Y,��<���b͔�j��LJ��t����}D)(�	�E�H��ɉ�և����s��<�$9�e.�pWX�����J�0���ꉟ�gr���ᵈ��R��`1KHZq|q�,���7�"*wC�r9�k���. ��r�=����l�r�sf�΍c�
��^SC�}(���|aB�� f;�&X��M��rS�]�\������mR^�a�t)���DJe���8���K@���F�CZ��S� �[�;���*f�K��g�M�
@�FB*�M�K�� �Nо��v��E��u��I&{��F������(ߨ�\)"�vM�8\S]��w�:v�bBm.1ʲ��r�8O�#k� ����b-�}��X	�Ƽ�/�I-�vV[��ݎE���ZT���5���s�!n�J� ��mwӘ$�7�!�i���r+t�'�o(�c�E�v��@�ؒ}� ����[�j�$�*���%Q{yx�� �ϤN�S� ���kɓ~9/���fZ=ϲ�J�cp�V(�U5C�F�4�-��ҨӢ��]�R<7���!dGï�sjfܱ������\��c�m��$J371�69��h��/G�f^dM�'>-��f�;�~���,�|����'��3<������P=���ћ�����K$0�&���K�v���3�9	�j3��^	�p�ߏA����vN���-��+ �z!1e�D��<����D����0�]�Iq*�ү6��UO��i^���rŤ�eN2<{�?����
�FJ�ip�T���?��9i���>���ת6�ax=�/M3���G5�;�p/gHd_���Zv�F
N���L£��0������h6���,Ab�$�%��V&Ep9���m�l�r���^"�iY2pb��a(�V�Z�;[PL���<�`4I��!P�u�D6�k	�sA���=�V�wMy,𜌺�WK����䂻��b��0w��1Y�9>��W[H�D�N ��1+|�ޤi+d�=�CB� IW`��'V�/v�B%3I������ U�����G^��X&��<��(c�(ٛ��x8���I�_b��xo�F��.�0p�k���)�T����Mϯ�WM �9�1�^
�W'U��=P���ll1���ʲK�K7'��8#�S;)�+�+�-��yI��e���RX:�Wk&�W(ݒᗻ���鞶��Ǽ��y��Ѓ��&�Pw�/a��k��Yۜ-� 7@5W���9@�D�k�eg�:��8i����!� 09�R�\W�lI/�L��!9�MV��U���&"�E�Y� ��赲;��gxl�(��&A��B���k�Ƕ��M���9:���ˬQy�I֥N��Ċ�!:��j��08/{��5=LCX���t����-��g����/����p�y�RT:R� �@�U)���s�/�9b�'��Ik0S���j5�d��N*a���II��N��X�iq���籼;�ф��VM��P��z?4*܆��lǺ��ǂ�3��'�yLv;�|C�4�W.�C~��n��A���s���%��m�huS��٣e�kEC�Q>a�2�e_���<#	���h��y^H���%{��⫓�X����r�\�%D�8ɹW�� .�L\�H������iF>�	��~=��fu�E�t���,�o#�/³ֶ�<��(�,�yG$������b��H��{<�:��d�������qz����S2�]4ϧW9�/���p�\���1�bv�O��&��Ʃ
ig�>料�+���#⛘�lM����:ӕ���^\��@֜�a����H��k�d3l7h��	�\���x�>���`@�Fx�Y�1�%=�H��ß��#b���749��e+xO:l>�� e�e�CE��E���US	*���l��S"��N��f4�)9���XP��e�fȆ�\�;T��ߵ���l�H� ��f �&��N3#��ler)7����5�s)�b��yR�m9�������m���YjV�r��<&`-���j_M��ۣic|:壿��@1���uM�1��щ��Q�ٴ�DT� ����$KAgd͌N�}��AY�~{�-�4g�ޕ�#+hIK⯼��2|�����{X&�� �t�����Ψ�bw?B]���i@�oP���JN�8I��'_��o���<U�X�K�]�L�wa	�Wl'KZڧ���H��\��9�s��c f����[̖��V�Y���s������Z���~�P~���&K?ph��@��-�Qؕ��l�i����u^�k�W�ٶ6_���E��XcF�`��;*��M������"Dk:~��J�������[jB��0u߶e��������v�b�B���@��z�~��BW��i/��m|p��=��F��*8�K��"s��rۺ�I�bu���*��,%6u�E�(K��rbUc �K�&�0�m5�NiT"O16���o�X�8�����b�p��Ձ>�e��ON5��̧�kzH�7bd����l�8'<_\{��T��^��Q_����eCԩE�%Z�����[�Y;H{6>C��H�Ƴ��M$�EAsɒ1>v E�-��A�������?�:F����)@�\L�#1�P���,!Z���@�]91���ˉ�|�������̒tV� T��O|���*z����:1E���Fn��>�?t�}��Cu ��J�j�G΁�[�Ϟ����W�byT��ɸ��a�(���n#�B���p��o,È�鰧�7��uX���jU�,��9E��kDOr�p3 =r3F$��¶)ssEH~���8�%D&B�� �$")�v��$�W[�`����u`b�Ô7��޶�&�n���V^���j6{�����'�e�G�$�w0���D.�Ѧ�~��q�m�.���7��J�ADF�	k���*��=��ʪ�wsm0�n�b�b���D�p"ͨ�1RbK��p��)�D��=�
�8��$hM��Y������
1��X���BW���_�}H�{�6���ӭ��[�s�ܬ'ӕt�\$��^��g��p4�p�����	�|�ei������%c��-�Zc�k��2s`�(���'�҆�ܿ#Z���3�K�b��*���6l
�~"xu�����T�e �k��-��Sɾ�hZ���g�g��2|��ͦ������Z(��tZ0f!l�'�0��0�7�!*�h�`�Ҋi�2����,�R�o!k^�V���O��pHb�%��D����:�ڎ�b�r���jY�%r�_,���	��'2aܝR�q����҃�ֈ%զi℩�:<���-v#�M�t
�\��;�I.��a�j�tǡ��p�m�v���b��͈	+�	0������,�T^o�Y	�ӷ6ua��������kAj�=�;����ի��w�����1=�����l�[:���R��a��אjw�'*�Vd���>mG  Yg��#�77<�[HՂ0UҰĊ�?O�:eg���-bݩ/�[kAJ[A��P�d�_���%#]��sQZIܰ���t�O�6�6c)U<�����J�r����"/Y㫫�A��If�\��Uk�4l��I_��ܚT��&�,���(��c6��glw�ͤ�+���ui!�L�� ���[���� ?aX��g��@�O�ٛ�}y@��ͧ���D
�E:E�o
����О&̈́��d4*�ZEA�K�K�Aӣa(G�#�-�4��Η��3feMj��TD:��V��q��1�=��� x����x�������!@G=�:L��$Bs�}>U=O��^��Zp2k�{��mh�����}�K�v�98��R��@�����4�8��|`7�?#4��S��lư=,f��el�y�]y�~y;W�A;�v�S�v��!(M�~��꺽^ݓgx(]E{��F �F�x��}#�g���a��P����-�3�^FH���s�����={�Â�7[i��|��A���V���BNV8�f}�F6~
-�k�x��I_��s��z�Y���E�q�5w``��W!`�[u��~�,���D%j1Ȣ�	�pn7�|��-�G�e^l�Z��Hi��)rn�G�R��qQߣ����hߘ�z�j�x��LT��=lH����I)/����{�Jʢ@�0?��EM�^����j�2KM�#՚��6g�2�ܪ�������,�ՙ��"+���S�+B�	�g�0}�[�ȓr ��ؼ��m�6$d65ˋ[�S�H{�@NZ֡��?�;���MR��D�*�ѷ��U��-�~��l�]'���g-�1M�[;%ض���q+V�&�nN 	�!�����s�ԓ�☠�M��x�f�����W�=���4����?�٣�WǥRu�N@�LV�η)��<��>�(~���u*�#�{&�s��OTa��W�Q�I�FTM����!����s�r
��l��N)�zL��`Y�sy�lF��i;�����N=ǟt�I��"d5ԋ�6я��N�AfB[o���^+�r<�$i��8�@�A7%�>��Q�%*[	8;�U�7Q^���a��O�a�'�-1`����Y�zpZ'}���#�W��}�׺,KP�d'�(�]+��!��(p�C-;fz�-��q�F䁀�! �(�R�a�t����F�$�W���B����
.���)Yş���a�LZy�݀�'K4auc2�'	������y��<g㟴��?O癘���y�l�_E�NR�s�a��3��Eq���m&i�ϱP����\s�l�)
�Ϸݼ�A����G}�*dA��4�ɸ�֚-�/���N<��JO��~���R��!`L��B.3�-ݴ����j1�����S���Ϻ��v7��T�1ޝ#a�:r�����V��fɀW��;�#Vh	�g��:��0���ܓ�����Q�!Ou.���?iOH��7�\c�� n�4t��l�C��O^��B2�SH�Ϸ�<F�
���]q�ױ���r_̇�R�,T��JҒ�1h����o?��r�?=l��G�=���;�B-�~�xx����g�#M���7�J����(EB���r���(d�	�F$��_D*kL��s��x�6�T?������B�9���u �ޥ��ci�w���~�9А�]�pc�W~~��tq�m#�gH"�s%:a}9�A|���7��D�W���I{A�NA.����M�y�`�o@~�#��s9w�ӆ��h���]޳����K���=�kuV[� ri&�S�
�1�U�W烌�g���S�S`�3ܤ��_���O�{\L�J�5�yl��c$��p��(���>d�d��߼
	]��	�"qj./΃���jBvqԾ�n�M�@���!�t@+�S��0=�Z��H}tM5���00�߈u3�a_O�$9|v 94�M�
� ���lW���}}T?��`Z�Rҽ�����|6K&�������� �9�+M8��E�(RU�f�?�?�_d���; �0�G@6�4��}����Gb�RE�7Sl�?1;Qģ.n;�J��:5G�u���A �Di�2Z���0@�t�g4�<H��B�u.mkM`�����ՌFN�����jЪ6F��,�p�j8�P=���70���Ֆ,�*Z:��[�{�����lЙ�*�L[�v�Nm�l���+����A�s*�*��z�p�r߸ ���3" !�Ҵ!���.�71W^~Y����i�@�s2A}��&e�'���ȃ<H�<0�s����q 5�^'��������p��U� n������U��d=��(���(R�
y��[QGN����9��ԋ2�9�Rܲ@������5 ;叄X:T�]A������EeE�r���4!�ZjszvÎ���TNj��蓃Pm�������<�eEd2���̐6إ��4EY�i�;�b�y9�QU��.D�7hG�z�8�
��K�j x��;�N��n;�|ҹ�>�N��bmp�����!� 	���Y�Wߔz)����� dR�`9�-����8�����ՍC�G����A��n��Ƈ��7��M �2 ���;:h�1��JIډ2N����w���������Nr�B� s�2aō����h�_fD���M�[$�."v8��A!�"��b( �݈ښ���-��Aݪ� ;�97�>N���DnX��/����������C}�_F4�cd��� ���+�?̒�~����[����\m�x=�����4L��:���I�l+Y�<I���N(B"�&|i5f /*�f�-o|��gy&��t���a��D�L�[�+�z�y�a`��`�������Hߖ�ξ�W�(eOj�Ӽ�U/�&I$@�jA`[Y��#oB����'ڋ9�)�D����)`о|65��ܒ�t�#�NsV$�^��ut�֕`E$r���i@c��Q� AI��Y��vzX�6��*��κP���;��xsS��G��m��C�#_�����ju9�����N��	�`��U̒k���v��3����}�G��Kr���{��2z���GGΉ�BOb���Z�b�J+_�~��E,�ԑꪭN������<C���WW<˷l�m��̓շw	.���Uf�c��������.=K��}���_z��TC^��+���4�l�f��WP��O4|"���{��x�z�PR���
��]��_cH�uVB�y��,�![R�I�R�����	�c��(���9�!�-�St�.zr�G!|�/��WCH���&"��{!�G+<�#�iG�jG�ԥ-?�m΀�͎>�ɻ��\�}m �m{ݳ�q�2yDO�%�6`����ZH.2_�F0%�j��@;����;zm`����ϯK�9M�tp����8�[Z�IA͡���-������]��>�i\Z����6�xW���O�oiz�.�&D��D���9�O�dd� f�-Nu��0Ck$-u��!�ߐ0[��Ͷ��՟��Q�3j��e�uE��>O�_��:Y��v7|��ֲ%pױ@q��t�P��b��h�B̠U�M��k�J}��7��ʀ�b�b�E����kFyV�0�<�ޖ����fMk4����o]�+L�Ѕ�hrL�.Kkr���^rC���"U��iD�R�%�Y�0��)�v�1����#O�L�����Ш�^|�� �kw�\R�g��>&�}
���ٿhN̅��S��l6���R^�$i�����4�k'�:�>,���^@���QB�m8�.1Z���[���4��Ee��`�fQ�)̍�`hShl�K�a!\}�f��<ʃ(>'�M/���$��:�}:����8f����b��.}�b��0��W�7���˗�o���)N�ۄ^H���w�^}���a���Ӕ�X�C5)ʓ}u"# <>��d}?�XL��>l=�5�_{��}��7��P����l�R��N��0%J{�8@qS��D�ז�H�)��T���m{S?�pє�d�5�/z��I�4���l�g��,A>�.ƊgK�D�A�js����	����>j*��u+1��@�W��ȕ���ͮnMP�h���o9��Lݥ���Ƞ�G��o~��>���z��wDq�G1r<�hI��3�M��[��)���bZ�)�Ȕ���\�u>�H�c c
t^�I4k�,%l������AHѳ���T�_	�5"���(�U��Dn�츗��*�v����;Q���#��Y�jYqh]�r�[���D>�#cP+�>�2�l�{>�u�/N�z�a��2�Q�x�L�#o���.d�V�@/��0L�,-��3��y�[`=��X����'>.K�դ��mbb�-�5�0��1?1�۞�&�&xx�_�䜼��٭F��j ����Jk1%�@�M&3S���d�.����D4�#�Su����!��dD��atZ���7F��(	�/D$(ko�ɳS��	�Yە�օ_��E�c6��a#�'	bK���&Km"w�3n��������y����v�Đ�l�C���
�H�ô[�ݤz�f6"�
%��Y��A��z�cf��I��U���7k	�ݿ�M�D�hpY��6!5���該s��z90�X
����%z�z�j�9��(��Tx,M�d�,�����	�u���HVh}��]��'��U��P�x馻r�]�,h���:�Gq�QDFA�i�#s��p�\1�^��M�{n�ᢅ0��� ���{Hq#d�s���w)�]G��Ѹ�7�y�s����sE������t��@7�hV���?s��Bv�ܗ4��}M�^X�ozxCR#��n>�A��'�^ ^T��d&ȐA�?��]���Pn7�qd��������\X1�f#����88�An�rY�_q��9捱h�7n=\���"�y�����Z�D�\��b��#�|}4�ip5�KY����H~y���|��V�v�&�Iw��޼O�K��{�I���-A	�g�
^�G�C`������.q�B<}�qe���P�z^
G��� ;�WD\�� �u]��	�� �%��`:�!��9�"lL�;��x)3;���.E�t�e@p����������OQq�>�iȋ׭٧ߏ�J!��z� �/+O&�P�yցY��72��Ӱ��^��s����"j�/��t�5%.k{�p��Z��O��R�Z'2׾�@�	�M
��Ewլ�2�dś.�����Sox�
m$!�b|$B=,.�s^�΅6RU��#�����Ip��k�7������w��KE&��Q=���6�k/���Y1�饽���_�y��$�쯑�k���r��*�&�(�v�'���'�hC��R�3�,,���}/�"��A
p��W32X&��KxZ>�7�Hz����Ҥ�$�f�XW���:^������"jR��W�Cv��(��Z��	�iF�W텓�4gH����E~~B�՝.�S�	�O�)MGm9� �s���ơ��n��$�������`Y�8OW:l"��ڡB��@�J3q��Ļ�o��?��[1N޶l�c������f����㋬7�j��F
�r��B�Ί�fĺ
>������ɃhD����;���l���zC<q%��'��u=uRK@<�뻓 �e��rѸ�m�����_�e&��2�NG�RvՍ�������t�D]�e��}\J�m�Y��sͅ
�f�y��F��`I������l ����'(��`k1U4%�>"��-�$[XV�#,�fK�E���(8*iu����*��n\��[���93V&
�+#�\�m;���p�la�<���iZ������@zbyW�|7��'�M��Jϥ3ܓ��gF��5Ź�p� ��2����aM��n��?��ܤ�p𸤔�{0@I��C��N7���#IY"0�����:��vDQn��<�N�,�O. ;�͖m�}�
U�W���+�Y����
[��⛮j���F�&;��jE�>\�=yy0�}�v�E���-��Dg5�ap���Z�d�G����� �mz3՘t���Tn��q�s�Ld�QMX���%�GNقT�y���
�|*�8����]��?�������o�~�I.��Pb9�ױ�.�9[�������"��0����5�<Y���i�l;#��]��NM�&�Ki����&�=��r3y̿�
��B����O�va�_�[���?����R��~�c6/�x��1��G�ĸ��A}�u]6�:��)ލDU�L���,�{��@M�g]����T��ٷ�w���&�zZK��7^Ƞ�����n�~��}�y� ����Ƶ����e��Ђ(�EѱbE�y��%Q-]{�v�N�=�n��v2��,YȖ̊U��"ٝ�Ž�B�2 �qa���s����yԩ���֦��)��������r￪窭����jȆ/�����Go��*缎2K'�N�B{��8��揃�-����dC�?������ �yF��P|0A0���sd�:��ߪ	����us0���IqL�Q���v��$�U����[H��
����jp�(�n$~v�6A{Ġ��n�j+�%=�J2��k��|7 w�3O�ĉҀx��0T���{T<Ԥ���RЭ��1f������~�%�[������xcZ��:�x��N���%U�g��t�a��S+��.7o�Cz�c�b��Yz��I���{*2r���R��e����P_3�$�uj�/�
�	�EQ����m]����d�t�����z �W�:���\\x���rZ�U{x���(-�%3��(��Q�,��ֲ�8�_~Y�W�M��3R�J��v?�Oh��&��~��Q�D>}�7��.�AI�n:R~[��}FxI�̰1�s��ӕ�i�rӱ�_�A�+0NK�+4�/d��F&�!�_����j���jR�}ˇ�R��r7V/�9�لq]�rWAE_����B7Ô4�D��5n&�cӪ�c��}�;2co�T�ջ~z=���#��� 1����y=?���]�J�,AH��@�աH�#	��z�`�e�4�M����v{}�Z�án4w%�Y�L�B�|��h�W8��s%RNu|Hhm��us� ��F�L���?�b�+q*�0�]�x����r�$�C��;C.��,���)5~�ż�x�[�d����.�p�9��e_ݣ	0M3�����Hr�2|�t��*.^kw�y7�J{%BkJ1R��x��6� $�_7�,��^ F&M����_��(���s��r�.��BT.$�񽲕^���%��K��4i�@��d�;�=e���q���'��ԸmH��8�@����8N#:��Y�3�=�UV�F���n;���ENo�h������T�� �@]��N����;�`ӵv���Ѡ�5z�k����ay�7"w�{h��DL�4�*��Z�3su��S*���gQ�9���x�����v���ϧo Љ��r�+��r�k���;�6<�ee��t+\�IN�6�.h��D��We�ۓ��v�a/
,~�T��o���m,���(���$��?�����nG9J��{a����|j�f���~*��o��{��O��*���@4��%���U�#lf&)�/�d̴���N��	#g�*ha
�n��${XuR1�A������ZT�V�Ug<Ft(��k�ذ�y*�(��\�{ܡU�!P ���(T|ʹM��p�X�&��F�����h�:E(Ah+����sX��"�%��*���V�^�� _�����=*uy��@��EÅh���w^��uU}�;���Ӟ��ʻu����L�U.�f&Vs���~���o����F�7�	�x����|��z��HFgGI^��~0�gBI�Zh�@���L5���]�=J��r�����X��n�s-�F]��n�n�I�T��8�fZ�}���9A���㑝5Y?~�a`
�rx
��U��7���e�ǄE���&k&h5�6Z�|�ͫ��!
b_K��W��
B�I�i��� qg%h�l1�]V��d����<���ݮ�RB�J�i��_�S5��y���ц�q���UҎ�(��������xs�ohE>l!C�Y9U�w��+��J��g�eP�"�H��Ň�>v3muw�ub�� �؎FK.��ND;�;ҷ`AK=��z2Ǟ�t>+:�W�+��2�|;L-�J�U��8�w#s@N�=�&�R���X��[���g�����3� !�t�U���_�Ema�_}cb�RL&َ�a��`` 5$ϫ�W/��cR��1gB�dm��"��ڧ$������v��(��N��bU��+G��� �Cp� ,x7���Y��!_Sc����-�f��@��C��B���v4�d�!�m8.s�l�>����XR��M�FȨ�Bs��˫���o`����+ُ�fA�>��rɻ�8cԻ�I��e_C���Z�� ����B2)�ȣa�	Z��Jy��U��0ZXz�V�-=��(Ķh��� �[%���?���w����߻�+����f���9:6�MWc!Qy�cm<Hڀݧ����[�G=J5�|2h*��E��m�Z�|O᧢�8O�Pee4
ʸO3U������147��\���a�c��e�
�%�