��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!��ߌ�6�u��S�`T
��E�E� -�5x8�ym�7�4�����Ƹ˲[�B�?�O�aq}A�_t�[J���J���z�KM��/��w"��ә^��O�4���n�����c�&J��Ϋ��	�z��-�\�Gs!���9��U��Rԣ�(d�k�Nd�L�4+�*C�l�Q|%�`��3gy�۳�,^�AsN�@rg����4��](���E	W��AȈ�Xu����/99>���[h��B���A����3_+�ƢG'���	<@�4��e�(�����]e����	��bj��0U�r'�s����*e�T�T!t�Dc��� �ୖ�Hq'���Xv�E�D�Y��~yN\�e�'�7�v5T:�h(�*�A�b7��d��=G3�)��m�f�iL��1�`��!���z�!�b��|6�2=]poV�q���:�J������|�0�5FM'���b!a�'�}�!]�n-��������{����9o�Hy��/@�:_�w"�F��cP8#�� ���.�i����������d���ۑ�:5o�<Fy}�����ڱ7�3��TI(�1%�b>��Wm�@����$dk59]0�J�/kf �^���V/�iz�+�<���>��|��;k�1EQ�e��O�޾�>�$�cD���qa�����@�(�6~�c�� �v�9�)��k*�c��Xպ7ia.��^��ׁńH��^��|4�K2f�_x��U���]e~֢P���\K �\�����7䐮�4.� 6oW��t����ͤB�h�}�ķ*j���gޛī%09\�p��	){��S�k��b_@"��8����O��hk����׭�����=��{����|a�l{6eYhp���hY����m���?��N� ��C��"�W�����Z�/ݐq�Ე�NSL��4[~s�suop3Ӣ[4���O#��j�JD�]^y�T�%~q[���VO����>S�ydm��Az'�]����?�����#��͚���u����9�J���� �E�)�<+�Q�f,�aD+x��5_�d�dBMA�m84��yk���^@�k���QO-�v������Vʴ!$A',���ހd�.�f5(��2�dGo^�ϒs�?�:!%T�y�`�S�$�^�s9X��\�ɪF0P%F��6��r�8ݤ�m�bt[��T�j�9�Ɲz|@��Z�ׅڤ���1�h�Z��I?%�T_H��|}'6����R�)Q�uJ�(�����}�җ�5��'�	��4~�6�A�/���ܿ��pMڍ#�!��R;pG�$� 2ͧ�%���Q��8Hv�Ϊ�6np��f�I��;��n�A.���e;����ڪ��"�ւ�}�B�����v�SI�_���{��+�KSK2y�o��q+p��˭�w�b�6�(���!��z��_�
K�|��l�k~MR� y3c�T��	��+�������f��1�7��VjzKɳ��mf��3��<���Q���"�����K�L�v����d�)����|�$������[�":���/^ßظ/�S.�l���ݡݫn�&����Ojs�F\�W��HE!�Db��o&NI+?[IH!�1�������0���"����Q,��VM@�ܝ(��	�7�:��#I��I�zZ2?���:�,�>zL����Y���5ҞN��Uׁ��>��Qz�0j<?��gk����=`���"��(����{mD]��&-���u�f�:�%�|����[WM��8�)j��&�N7@n��/9�dyI�'�S1:�E�`7�}�f�>\��sx��Z�F��������8��p�^�[*��|�s���	:欚���F�a)��(}J�y�ˬ�%�r�+�玿H�Y8L3��a����Q�t���l�k����<z��%��{b�r�8f<z��������h"W����iSR���h����O��r�z���PH��:�׈�9(Uz|��S�,n�B�M.�I;@UA&��w�F�]ˡ��W�3�s�~��|P<?G��jM��J{�ι��ݺ�$�?ގC�_�EQ�'�G\���g��0�~�o�����cM�J*ޡ���-ؙ�n�I�]!/5m�}}O/��p.ӏ��H���2xr��o<ć�������c�r	����7\ng|��y���6R�A`B-n�w���ķ�\�-��v{��Y�(��� ��;_�P�#:���L +��p@���w�!�.�XD����K|�~���'�m�R�b�[���8�^��g�i��qU�l�\���Cמ�D[!��y��J�j��r���X�3���<��Y��*	� ���`�u���|A�5�M5�~Ti��8\�G?\��
v"'�k�NQ���lʊ�����,(	�`�+�%�?fۧp�����>+p�,�� �@|�r�� ։��+s����m���0�ܯ�KTS�kG� {('r[��Lv贱B�m��5yz6Z�"��\.	�.��D�C��B��}}����7��]ŷ�VW���3���?�]4��A��Ҥ�</�p�:s��R�J���Դ�<5������������Ɛ��8����	;����M�<B91�y�׃'0�� 5N7�؊�j�5lb���[y��~�
��f���[�������g��&{��썕���\��aKb��-�HЫ)�qԐP݇�T���J�&�Q�<H1
�I���N���/�cNA��0~�)J'\	8fx���-�Ҁm/Fp�b�
���2�M7!�T����cї�K����L�醉G��I)���z�X�2�~z?'	��bm�!�<���L�K�G���4�$���k�����~�)��~��c���[���:Y��s�]� �7�B�_��ǯ Uh Y�0g5������bs?c���SY��5@�1��{�?2��t�que�)��ވƙt}x���J�9t�x6��(��v��˱�9p-�_3k���]I�⼽+"�L_�ۀ0��ɫ'�c�1�3��L��lO�yul��y��w ) ��f;a׳�Mhކ?j�$��Wq�2�Xykms��U��ۼa����� �KE�܊�oaz�ѯY��ۭP^���q���6��[AU����C���d�f;ߘ<dH鹵�c�+���$Q�n�S�0�1�$'�����8,-�b�~�H*�-M*�xv�M����=f	���M���T�2�ΈZ�煖:��
~���c����̡̈~��X4S����^�l�pyy��ŐNa�ßU]=���Ls��swp����8��Z�qԭ�,C��+�9:<��;���fW�n�À�j�9{Y�1?��8�����/��u.���D��G�rfmuy,l��AF��<W�>̘ې(%e�<gȄ�2��@�>`9>�T/��ԇ��p��Ą�>'K���R�$r��~n��g�x@Ω��WOB�mOkHT�,"�K�/65n$���k�:��+U���r>C�z���\4�(�e�7X������W�bՐ�|�@C&8#��v2�jZʍŝ�Ѣ���J��)�_��i@Z<zq$ač�`��K��@u,�Fx����g`���#�C1p�t ��z�@f@����R_q�~��k���dzc v��M�������E�O]D�� �;�KD
>w����l-���[(�`Q�<����� @�vK���+Y�K�(��:M+�#���yw~�>�g�d-F?D�NO
4;'Q�iRܫ:z,�J.�ϱ�[.j� ܤm@N�@%սN�Z�B
�+��Y͉�^�T���10Bb↦�60.e���,��,��o�3���i�:܌��k=z����Kc��N�9f:�k{���c�Bxi8FR�+�ǽ#i��4@� F/n*I�Qmh"�BH�yTML,�����]I�y>8#�X=b���H�����h]������2�*�M��]���k8���j�XQ�	_zj��q�ڃ����y"�93z��@)eZ�v:�����N�vʀ��8[������ӆ����͕#'E�!�EP���:L߾7�kF���{�L\�o�y>��"����Z]|��2��������)h�9=2 �Z��#�������k�K��hu���XP�8�7�����̰_�ڙp��%]��͇ts\ɫ&�ѻr#1*��+�b��Ͽ(�[5���ĳw���0>I�7t!=�gG��� 'YJ3��ỗ��-��hs�C���k-���c����G(�+�40�u��Bo�Շ<h����gn�F�QiM�:�i	�<8��D�Dr[o����)��l(�jӞǏ���=��\�_F���+�u2X�!E���_w�!G�G"�W���|�����a;���6�/b����4�Q`�=o�6٪�.�W�l�ˉ��l5r 	��x����9o�HД��Wƈ�
��N9K���U��A�k��"�=�qrm�09V�E�~W��i���t>�ǌ���z��c�����>�G�0Ӱ�<zK��}�3�fw����G%bY�D�"��1mhL���[�¨��:��9:�n�B�b]��C�}�d�K��b��ѿ�h\�k�K8oQ�`~f����9��!\���}��n�G������ ���r�]���KkcG#��as�MO�ʁ�3b��"W�i��!�>Y���*�dS�$&3[�ĎA*�L��ҕ��{Fxt��K��"��8�9�@�S@��4}>�f}�=��*�]*1�68,AI�D�b�#�^�A]�̛����i�e���?lŲI{B��M��B����Um�m��Ώ�,D�U�Ɉ�2UMг@3RS�X�x%�Z��;fy���_ԤZ[LrB���,'S�	c�Q�Fԥ�<Oƶ#Dә֯O �'}2HiL�Ƽg���H���B����Awu��fXIk�;}X���(��I+�K�m5�����<�饃�����N�b,�2+��;�+�v�����lA+au}�G�`!뮍��cn��v��� 4��p���Oǉ�����,%㤴1Հ��,n�e�hTU�oLBm�y�nzG&��7��䟙k���U}.�郧��a(��!�\��(L�Y�J�����g�mF�3?tq�Z��>�;��;�[�#F=Jh���~$:I��q��roJ�]�&/���{��r�dݯ����.�k�q;F=����`OP-b4.�c̺�4�	X��o6Jd��U�OX(|��|˚�*��;|nb�_Eu%z�3.���;d�Z�a#E>���>���rB�?���jQ.X`�E���V�6�N6��Ԛ��~�W�c$����/֍��x.P#����K&;��('LC/�#8k��!6�{#M���|Lr�U��PJEϘ-���%�n�d��:upC	y`@���K�:��64�)�u��,��r�y���a���H�{�(x~b.����v��1�lɒl"�`(c��f�ә.f'������w�#ݞ��w��V�3͊�p*]
Ҽ.�.-�[aa�6�/�,�j9�zP��I���������%�tma���i����ه�L�=x�]�<��õk�� ��e: 9�I���׼#�����+oֻs�I���~���
ĨoD�O����>�tЛ�'t�T�^	Eq:��@��c*���P6����O|$��^TT@C������8��^�×rI��b�D���Ʃ���]���P��սv��We�r��>��4�^���ͽ���~�h繠�D �>�`{.���_���޾E�`)&�vw�1�7i��n�V���N��{��N�L1���ַP�#�8L�zV���k�'���1gC�*9l��D�D�����&�e?m��੧�EIG��ٹ�|�!7F������0�GV�ktM�Nwm��q��my�U��b���%&�יo��j�x��� ���D��&��k�u�90�4:���.�7��Gٙ[8��Z�u�����,Z�k����.��x�q��������Ջ�#4-8�=�5Ė��n�"ȑ4d:�lU虣��� �ꐦ���E��7h���#@�Xt��L����o��g�oї����DͰ���^�Xp]$Oz�M�	�"��~��3� ��W�����'����Y�lh0��k6��~^�����B�> ��,���f�_?�S=���ɠ qf���h�#E��q�./,��Aq��H������Y�]��""�[��'q�&;z1���̊��L���sS�,��<f���%�/��@��5�vs�a���P6&mfZ��GC�x?�_��ܾec�"��m�F�g舴�e������z�����H��X��cٜ!�ljo��;Z1 ���=n����ɫ�h���Z �gي�xfX@x/�#�����Wur6W_]��yw�'}Y��\���K�Z7����2�	��,[��C�c �de�C{��4�6z�ZrEY�i}d8Qм&����c�[��^^�1�j���d�ɹ) \��4?���	�Dʬw5�d����X���N�}��t���"R���:cʭ���چ7�|�Kz�ck7���|c��e-�j��x���p�+�� �i��5
���4}ҹ<p�rc�KV��銛�?4,�>�g�`��r��}�u$k����b/Oܳb4���KЙN�C�;´��&~pR��z�'�X�'��\�b�?�C;��6�e��<	@��J�U�k|1mX�-���ę�6 �]%J��va�'��0��������5��q6o:Y��X%�:V����X�OM%�~�&�G$�@��7ރh�r�'����qoR����	;��T.ɔ���u�h���yZe�tr���4~W��Kr����9`VR5p�q�B[���#'�q�v�s^�U�nr�k�ϹM���ݼ�Zc�g�V��:�0���{��-�E�.��Ě>& 11j�ٻ��|�l���13������U	��IC�28�K�	� P�t�v+_C�]B�oI�od��<v�IId�7o�٨hZx���	� � �<�r���qx�*/�ګ+7h��n���!�j�w���D��Jߡ�ζ�+,�]  L�nw�Wl1����:���p�1�ɯ�9"o��'?�W��з*-����G0�B`�=����/���9�[�AS�^�����4�8F0t!W��"sA�H�lZ�)��ix�5�7��+�t)J&d��ׯӊ�lF��E�Kve����@0��Y;*'���I�X!���%[�L!��Q�X����Z��%bB�4�G�zA�hՠoYq��Eij�����l�:��W	��ȏnZ$��O��p�L��z.j| �A��u�f�Y�`(��l�����AG�~%:�QJ�e�:��5������Y&<��$����~h&����^e�	��@���)��l�
,�%� ��~��V��H�ň:��ݑ4�<�A�%���^�ȗ`����6	�Ā���]�� �i��\�X�r�(I��I��ewpD�������-��\٣ڞ��4�:Ӻӝ���an{&za�FΊ8������(�#�uz��^�?p�{�*1v�W.��"���1����s8X�G�"�9d�dޥ�5��z')T.7�.CT��t�|<kfBS��ߋ���KGx����G��ɀU��5}�7n�r�=Y�΁q�`�2�MM��oK#�K,o��z�u�����k��j�.�/���~�YmJ������xh�q$�w\����w� ��_�R�HR0�����<��gX���q�86^L�U6I��# ��U3/��$�
������fZ�#2k܁�i�Bƃ���R�%������� w_�.�@~rX ΀8b�J#YQޢ�P7}���������m�3����׹��:�|G2&�3u� �>�z|��O��ˮ��qp; �́{��\yX�ҨyMaӾ�ոP"E�ޚ�\r�@!�6��%���/V�n�y��H�bp!�H�L��}�Y�t�'��<�rOI�1����d���l��&N~�6�ۊ,_ '��ϯ�$�Y�
;	5���0E����W�V�2c���Hi��S2iCn�̔��(m���a��z�X�F���EQW�Fߘ�d����A���ӤV,��j���!D58r5�[ƿ+ai�ƍ
��o�Ns\�#dI1J>t*��XW�4N�����/v���q����'�J��҇�=�eNł�a��7�f��g2���M�B)hё-B�+*��h�e]�_Y_��������zV��pL�X��ݼíJ*G"r'���'��%t�����Eݜ.�Q!%<��=��E�B(�u��Y���R���k��K�N����~$��>G^mYۨ~lZ��r��?�;�dn�Տ���hH�!�L`���eD�U���[���2cQ6�c�JT��6�N�v��#���נ4~1������GL���W��O�V؁�گ�P���3r*��/G��y�qJ����:��I�۰׽�x\Ӟb�*��+}@=�\|-����ъ�J*�[���<o�iߤ�e�|�+�Jm�\��3�m84��g3��b�瀐x��aIꂪ-�b����{M4�
���8.D�A��`t�$=[ס5�L~iH��!~�R[��(.����Y.���4	+�iBz�5���ٸb�8]e'�D�#C(|���-���'���b���{�:�Zۈ4�6�ot	�*d$�]f_�]�\��*U?���(����v�i�EToWB�&Y9j�\�蟊f3)Wd����4����u���y@3�`��C��#ln���i�K��`vp��ՕR]���ȃ:�E�1��H<~F��v3O"נ�Au��8#F2�?���3E��1�VAm"�5T]�I����~�+������N��1\7����h�Qe�jO'�T��'m�S�4�͌[m5�H����P�ٻ_�=��[}�d��1��%��۠��,�w'�X�RwȂ	)��+����;W�Q�׫�1�	P\��MDMnM�jH��7<���X�K�֤��wջ���|�q�w�ޓ��8��u���b�/�s,�c#_��cpԣ��l�ݥ���\#�[R�h� ��$�?�<�b�fB\7g�M¼�����
mѦE/�|�V�=M�J��}�{�U?ET���xE�C�W��4�'7���EJ}���8�3��Mj5�_Pq�MJ� �b���}f����� �J�C�s�߮�����g�GId�&���փ�e����F���l���K���Q�����8����?E��)Iv�x`���}���$���.n��F�y�� ��� �b��U1Q��l�*B�����(k���D���/����`��\��4�MyVD�����#�$��ּ�'�q �!@�=���C<S��DJ�6p�L�N]����޿��?��ڟM�o����RxVE�Ø+��9ry [#�	��*w����@��g�/ �-	D�*u����'/�H����
���Ȋ�%���~~=$�I/�1�v����U=�=(@u
�Ӥ�/�Y���H�`8ݓ�|B��eS����L��1f�
���H+������T:�^�^�Ԟ���mh���
�����5����=�<SK]��9p�2����B�`����������HH�#� o1t���qC^�M���u��a��^���Kr���düx92� Jr|e�T}���EdE!�u�G(P)���XI8�v@숇�j��yW��7�f�޿�ЮE��G^��@���f:5�{N[��T0�W�\�k��G���;�Z���=�+��Wɖ�����>PH����9�l���fq�Q���7�R�� f�e���7�=�B͖��R��w�#��ۤ�3=am�g���b��/{��+9�Ý���6�j��w��:]�9f8�ү��hh��9��6���`��b2W��@��8�v���K��ڳ)%���J����FY���^��q�&��m�uA��v����?"��CBs�QG�U�[�;�x�$��̭^�[T���&)D���x+K�J��.ɀ�k��Ft�c�ȫ�
x��J�[��~��H~���ɭ]��c��Ob�æ�[��Z���Kw���t�I��UQ^�@6�sb�w+��	�%��bT���p�F��?�'�/�l�7@O�X���uKO3+MC��+��_�G?�J�SLΑ�=��|�˂�5�x�)��+$�dǬ��%��Y���1['�>u屢����Z��ZN�#�f��Gl�YU?ob�O@D��q�6�	F6B��l�O���Ī3����4��AҫυKJ��p%���22��U�|��!�p[���ͰW>��l��?�9o����( J��-82/���&BHTP��`44>�����`��3kf����U:��xC���������(M��� �����9��/$]����X�[��͙��=}��5��@F׋�֜�;�\4�/�a��M�,Q�7����<�= `��`�ݶ%���%PP%E�:�e��`�`v��Z���:ʮͱ� �dR+Ù�=
��n�{&�C޻��5�-����,�`��^��P�jD��|�i/����oH��g� �h)��� ��X&�����A��޶/�Wn�Ą�[��hj?p��0C�/�� �|�מo�Q;n��i�6�\8�H��X:^?�pQy�Q�ڛ�6�{���K��ŏA�,+h<�xl��� ��,c�X�+Aa�Ce{��K�
Šz�dt��U�e@�n"ho��;W~�t�*��[�.I;���tO##�XH4W,���+�@����Km[�"��q
GS/R2�DP�0���k��C�:MWB�>ɇ_�����0�D�Lv	t�>zWa4���a�b1�BY��r����h�����R�~��9e8*r�=�#�X9P��j��	2"Yf)/ 늩���$���!.�)QoI=2Fr�)�7�XЫtqӴDi��������qGq��V�K��k߬��H8?�WQ�A���졹�1�c�5'K!�:�́N,~0c�P������H���= 2���K��`�撙B`�f�Dӱޒ␢��{!�ǋ��)H fp�(?h_W��A�:^<�oM-�PE:�m�1B��L�ˍ2��U1CE�R�U��MYĭJ�����
N��6c�(������K_M �M�<\�q�`c�E���~�(5���Í�.�딯h�׌��oz�Nd]�;T6�5�ūP� YP���[u-rYZ(���5��������+�j�#��<�~6����⵵%`�O3x( 1t�"�򈭛�ӛ3�*�l�,E���#R�T��	�:,��q��t7iǨ\v�e����b���5$�������b�͗�k��l�wեpe�0yW��������\�,�vHƱ�$x�SIe�wq%�
�5�>W�~�f*@�Rg��Z]�>�1���ℸ�d`Ta�Ѷ�����ks_��ՕU9s���##�?-�7�x����Z��� i�"�0�C��*�sJb�@s��	l�z�Efz�������6O��Dl�c��C�CW����9+��կ�2� ��I������ �3�Վ�Y����4��ƍ�B�%ț�g�3�U�ւٍ��A�^�n%�:E��)6�Ui��a"Wz�`FGq���h�v��١����c�h�7��ϡ�/����E������%�
B��C�(͵e)�t�0Ә�*k�rev�����0aS�X�3ٿy��?\9�?~��Ak`�ND�l�[ŁS�(�.������Y���E�^�/
����C�`���ңA��b�!�lq�˶*�������69)�z��{����ڞ�,b\F:���o�2r��`��:T�!�{F���$O9�@�
�/���Dc�w��P�4h���#^owD�*���<�6���f�gB�U���㻚� �$����]'�y��k�A�|*2�1��Y��p��[( A�{K��av|���c.]�� ��H�V�w�w�m�(%�g�2 Qڊ����@Į�J�ΥB�BlC�B ݔ�D��@G]��G����9X+]�?zON��j�n��F7'�9�v@+�\8�m83�4u>���ܨ�ы���:ǅ�����Ь�$����Ă��4��I�uk�$&|�4z�,������q��A:���-jK����B1{��?B�QJ�uᤩ>R��'(�O�i(��9Q��w��y�e7�^c�]r'\���4b���#�^$�ɺ>~��q>QJYR	U�Qj^ī���<Ǒv,>x$���bEڭ�!��V��%���og�L�%��?Q} Y�I��I�j?�8�=`	�����?�\��`!w��\�Ο���
�Q�d��)Q�Y�6�$q$��P;ڨ�W�ñ`��� T�u�D���֟��r#�Q��U�rDC�Y�, ����x�J�u��EF�\����2�幹��/�J	*�M�S�P�) ��ݰфP������LI�!��:?�F�duHzS��Z��z	��U���~0@����ێY�~y�S�|Q.���MPN|����df�E��g�t�/:��W�	�u�T{���,l�o�F,t�,c��Y��\��m[�Z���Fi�ZR��$��!�:I��jnûo�8YpMI�I\nT��89)��sEd�󺦅&l_�]b��_i�8��3pZ'�A6��b����J�,V`DMG��~�\C��S#�AN1��i�! �|2��p0g#$���~�ɺmYz04��S�j�h����K ���?��Z�/v;����~
�YC�b����%����&b�r�~^�����|5*!�|����}��O%��J��|��mScxܻ�J�,��Z�d���\��e����2�ۙ��0P���<��t�=%��+��H���D޸�}�޾3v(��A��my�î`us�����C���0��n�	L��"�wgS-���޶S]0	3D]scL)H%hЏ���Gm���t���Ӵ�UZ�ԚW�#���T�,�b�=�	.��M�8>�0�����ɬ�Ɛ֝/+;G$O����f���=�{�׻{p'��ȴ�6d����'�o�!x|AI� O�˸���i��2N�cN#�Q��9�S5/[d�:@$����n�ch@�$$�M�q�^`�@��R�s_�/��PQ}*�?tX��]d�-s�?��zy��x�P/�
[����k�5S�B��'���Dz��ʌ��A1IHqL.����uO*I@Xӓ`>ժ�6.�Ӯԓ��ww{_�V�/[DՁx�j�@Q;�$o�l���J\bj�7����ir%���X�A����N˘���B��v͋#��:�*���/�8��l���G�<C�FcE�� ��q�����Y��SA�H���/�ݨ>��w��[����r+G_ڥ�+$�z���:�J�F���OҊ��(�(&��/�O���6+���o���uB��c��Z����G��l�O��O�Ҳ��mǖ`������)��ʇl�(�l߹������]�&D�7?r%�M0�6��	1or�6С��u͇B��vK�Ը� ��H��-Թ,ae��m;��D�.f�z��xϭ�1�L���[_�j4y���K�e�����G.S��j��{u���j��*n�T�w�[!����c_RPy��~K'�u�n�F�����_�{��t���:�Gn{�\n�����H�P��#���x;���u3��a]�y�<��(B �K�@W�� q@�6R�@b]�1��b�>����8c�L��z��1�����)����ϳTF޳�ň�~TRR�mxY�Jm���y��M�ZKT��S���!���r��ֿa3����c�YgR��-��T��"졬2�*~ n� Cꁃ��D:�ڱA��Z���[^\�6�ND�KEb�q�)r��~R������䙰�>6Dg�*�#�Bu.Y��H ����o�Y�~����#j=��͐n�X��gq<���s]��(gT�K�d�%v��DQZ�Bw���nV��B`�eEy�CA(TH��Y:TY�������k��T�ƫ^��XIC��m�&�N�� ��������O}�p���i�ᇏol����8]n��1��l�l��/8��]���g�����@	*��ȓU���0}<�зƂ,�g�a�1�)��3���4���5:�T#���y"�R?���ǌ��Х�;"��i�ڱ�*_�M,ɕ=�)�b&n��4�����P��O8���P}P�'�0#�L
W���_f*�k�uw,�!0"{Iq��u�˵U�T�q��g�z��e�b�� �E��˜��1����[���Z'N³���'1���z��j��
r��Y��uu��'�4=E�
-�Ƶ߰JE�%}�)�+�bL.K �l��
�3��S�����Uz�[1Oo�>!����:}iǿ���+�P:�0�,(�jk�����F�4�x���R�5�H�
�x�w��5�2�c�^��5��B�m	&�P���u��H�X]�o�mJ�����{q� �m�oc� O*�� ����^*7WO������I,}M�X���av�o��Xѣ�%���*y���V�%��������,��4�䤰h
%�������j���.���򳝐[��z�Z;M=�}��
XU��U���v�N�$��~��Y29}W 5�0¨��h$f%��}��K#�w��d����
�pJE[UZ�&�0������\���ȕ��� s�0�|}f�3�w�Ӕht�<j��=f0`Tހ�ߏ>�:� ��X
���qw��xAU/&-�j7s���_������YFd5M��?��m�|蠛���{0>r�$5�|�*��M�����-�{�TV*!���1ZL�!�Y�ʻ*�S���K�1�4�'��5|�a�a�G�[;���*���HbܧڷG�Xg���K�D&��z��E]��"��t�v��>�5��|�6j`������c���fG1F���i�8�m�e�;��0\�)���ˊ*����,L.ߧ�E��#��D�sR�G��R�r>���J��S@����
iG`>Ju�X�ʺ��[Yot�I�����~������oG\3���fh��YRzAEA���
 �eʱ6�q�lC,wz�E9��O����o�6�,��f����9��+xUO>Ͻ����<n(�@9��n���m�����F�a"�
�_�*�+�J�$����:M�UV�	HA@p	@M�_EJ"��î�>��6�H�L�_�U:��C�L'Ձf��1�zhX,���z�\U�"�=�4J�z`���<ٳ3�d[ UOgAА�m$[0��Z&e�왶�r�$,��;]�I���	js_OBY�R�	�:�Q+��#^�!�s�����A�w��H��ҥ��������N=%!}����r)�9�ɲt��!��	)
�n`~����.>H�sr$�Z�����*�J�&��)i���K�ׯ��d{,C����#J���P��=@��պ,��>��\	��ߑԬ�.��o+k�LPŌF2�a�\�y=����mB�#P���g���ӳ4"{w!6������˂���q���U$�����0���x��nL��e2�S��C�{�Q:?&?.1+�x�M���0�`Q�Y���2�s�+T'��p��<�����w������"����(k�\�K��[���>����k�h���;t
=�����sNs酸��� �^��\$��a1*?	YӈP@��kղ�q��"x�3drH����Qi�g�[��DVi<^�r �I�!ci(�a�0i�G����9M*�Jtt?�ݞU)�)Su��-�Rvr. ��,�����0>�f�|��������X,4jґ�4�ѰZPw ���/��y����p!�5O�j�g��<A�
y������K����g��7
���d�#h5�zyD�0��#�P3�G�-�a]ms�b��I�?��)�:����	`
���D��b)��sP��M�s��O����FY� ��B������<�*�����mG�ta'(l�`�:�K����Gg�EY�6��� "���]8�Z殡��lu�d��zgXK�@Nvw���)�M��pOkkf�K�b(�)â��
(�./��<�*��Y��ߢ�o�_��	A�a�6�
I;𘇤�ha�1Q	`�SSf
�Z�՞��~�OC:l0�fG�3��b����4�V6�bŋz �wv=�\n��5.�%��q����
{�B��"���G��i5�"id���ϯ��*�{׮�L&@"X���M���Y��v8��os�ܗ0�_ `�?�C��d���"~ށ��M�MI �!�V�����G��b�D�I��B��.��_�`	��m��Yh��c9'j�3��0��N�x�ֵ�e��R'��U+���(��י"Lon�DGJ�t �.��a�Q5&��F�'k'�W/H��^��X�BGz�$V�L��Xq�؀�[f����$Ӯ��>�v�֝�.iJz�>`�U�	15J��F�%�� `����l-XQ�	Ey�}��ś�2���m�{Y��0�c&Dꪨ�׺�6�'1\-��jqx����m0�ȥ�<��L�bV*��1��y��
倷�w��q�&�^M�˷�#_�r6�*0&� {������Æw�e�����x:��58�H�g��{|�V�GT=����f��5�̈.��-�	[(��J��X���&�^��z��j���-���2���L�ڸ]k?}1�-��piQj
0�U4�Xf�U ��eh�$�N?��X�� �1�`�����=UĲ3Ѐ�8���r�E�'v�Q�k:]"�b.�!!W�Ʊs���U�D�3����/<,�Ƕ�g��3��-�.�o��c�uNQ��W8=H��r{[�?�����Z:3���?6Ն���Oxd���j j��Ip�+�å�1n��L�GŻ�|�HgQ���K� ɥ���0މ��.E{D�T߂�Eҽ]�/�;��Ɠd�t�$�mh�QV�P�F�l�����i`��q/05f�ȣ�ts�#|*�MY��������~�-�v���/�1��AZh�vF+$`�@ŧ����_���y)؎?B���j���&C��:r���Ǌ����i��ő�k�t�� ��I���Kl�� t{:�����Fꋄ����(Z�\����4�z����	}.�°3��b� ��>�اW̆�z��BZ�����w�ۏ��{�}7BS��˶�z���K�rQ9߿or`%�M���E�}�vO"m#n���e}�F'�����bR���T�$:VK��ұ�@��l)��_&�H�`�G�(�&KcxrC��zx��g�^���܄�s��:�B�\�Y_���?��:�s����} �3��O�b��v:�b';�X����h��s�C����V�>�%�����8?:t [vZ���o�i'��^�~Ԝ9�	He�f����7u��M�BZb��iE�2*]��Z�*%	��/��V�ס��kiI1��jI��s;At�T�Q�ˋ!��h�ѧ�rZ�C����C�H��F����;���~
(M��3�*�B��ޏ��G��Q�^��6�V$����C�v�$jXggslQ�ة�vz����a�����n��߷F��M��f?�+����aG}赐����yp&f Zh�8�q0�:�L���"wL}&�3�yZ�l��L�U�VR�����\���VuX/�Ӂ,���/����3�@�PU����?�G_�3YQ�bÕ	LZ��/��S*;��xN+:"oGJ���b�oGV{���B��θ����Y��a=D��2�R�m0F�.��@�,x�S��pxā{c�PY�l��ԔA�0)��~�r�k�V�D�Zi>���$�4C��S`޿;$�!!di��U�h�h����;�OBE��L[Ҡ�Z�PrR����O|��c�̏|�誄�w�t��k�U�Ƒ'�X�����l)I�����\@��`?��s�W�K��Ƌ~X�<I��&��iA�~�������J���K��%�I~G�o�(,C��z=NY |�A��l�����S;@��4����z̧��� t�T��P�7."l���fOi����C��g�To}