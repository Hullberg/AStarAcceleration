-- megafunction wizard: %Stratix V Hard IP for PCI Express v13.1%
-- GENERATION: XML
-- pcie_SV_hard_ip.vhd

-- Generated using ACDS version 13.1 162 at 2013.11.08.15:31:05

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pcie_SV_hard_ip is
	generic (
		GEN_RATE : string := "Gen2 (5.0 Gbps)";
		MS_CYCLE_COUNT : integer := 248500;
		DEVICE_ID : integer := 4);
	port (
		npor               : in  std_logic                      := '0';             --               npor.npor
		pin_perst          : in  std_logic                      := '0';             --                   .pin_perst
		lmi_addr           : in  std_logic_vector(11 downto 0)  := (others => '0'); --                lmi.lmi_addr
		lmi_din            : in  std_logic_vector(31 downto 0)  := (others => '0'); --                   .lmi_din
		lmi_rden           : in  std_logic                      := '0';             --                   .lmi_rden
		lmi_wren           : in  std_logic                      := '0';             --                   .lmi_wren
		lmi_ack            : out std_logic;                                         --                   .lmi_ack
		lmi_dout           : out std_logic_vector(31 downto 0);                     --                   .lmi_dout
		hpg_ctrler         : in  std_logic_vector(4 downto 0)   := (others => '0'); --          config_tl.hpg_ctrler
		tl_cfg_add         : out std_logic_vector(3 downto 0);                      --                   .tl_cfg_add
		tl_cfg_ctl         : out std_logic_vector(31 downto 0);                     --                   .tl_cfg_ctl
		tl_cfg_sts         : out std_logic_vector(52 downto 0);                     --                   .tl_cfg_sts
		cpl_err            : in  std_logic_vector(6 downto 0)   := (others => '0'); --                   .cpl_err
		cpl_pending        : in  std_logic                      := '0';             --                   .cpl_pending
		pm_auxpwr          : in  std_logic                      := '0';             --         power_mngt.pm_auxpwr
		pm_data            : in  std_logic_vector(9 downto 0)   := (others => '0'); --                   .pm_data
		pme_to_cr          : in  std_logic                      := '0';             --                   .pme_to_cr
		pm_event           : in  std_logic                      := '0';             --                   .pm_event
		pme_to_sr          : out std_logic;                                         --                   .pme_to_sr
		rx_st_sop          : out std_logic_vector(0 downto 0);                      --              rx_st.startofpacket
		rx_st_eop          : out std_logic_vector(0 downto 0);                      --                   .endofpacket
		rx_st_err          : out std_logic_vector(0 downto 0);                      --                   .error
		rx_st_valid        : out std_logic_vector(0 downto 0);                      --                   .valid
		rx_st_empty        : out std_logic_vector(1 downto 0);                      --                   .empty
		rx_st_ready        : in  std_logic                      := '0';             --                   .ready
		rx_st_data         : out std_logic_vector(127 downto 0);                    --                   .data
		rx_st_bar          : out std_logic_vector(7 downto 0);                      --          rx_bar_be.rx_st_bar
		rx_st_mask         : in  std_logic                      := '0';             --                   .rx_st_mask
		tx_st_sop          : in  std_logic_vector(0 downto 0)   := (others => '0'); --              tx_st.startofpacket
		tx_st_eop          : in  std_logic_vector(0 downto 0)   := (others => '0'); --                   .endofpacket
		tx_st_err          : in  std_logic_vector(0 downto 0)   := (others => '0'); --                   .error
		tx_st_valid        : in  std_logic_vector(0 downto 0)   := (others => '0'); --                   .valid
		tx_st_empty        : in  std_logic_vector(1 downto 0)   := (others => '0'); --                   .empty
		tx_st_ready        : out std_logic;                                         --                   .ready
		tx_st_data         : in  std_logic_vector(127 downto 0) := (others => '0'); --                   .data
		tx_cred_datafccp   : out std_logic_vector(11 downto 0);                     --            tx_cred.tx_cred_datafccp
		tx_cred_datafcnp   : out std_logic_vector(11 downto 0);                     --                   .tx_cred_datafcnp
		tx_cred_datafcp    : out std_logic_vector(11 downto 0);                     --                   .tx_cred_datafcp
		tx_cred_fchipcons  : out std_logic_vector(5 downto 0);                      --                   .tx_cred_fchipcons
		tx_cred_fcinfinite : out std_logic_vector(5 downto 0);                      --                   .tx_cred_fcinfinite
		tx_cred_hdrfccp    : out std_logic_vector(7 downto 0);                      --                   .tx_cred_hdrfccp
		tx_cred_hdrfcnp    : out std_logic_vector(7 downto 0);                      --                   .tx_cred_hdrfcnp
		tx_cred_hdrfcp     : out std_logic_vector(7 downto 0);                      --                   .tx_cred_hdrfcp
		pld_clk            : in  std_logic                      := '0';             --            pld_clk.clk
		coreclkout_hip     : out std_logic;                                         --     coreclkout_hip.clk
		refclk             : in  std_logic                      := '0';             --             refclk.clk
		reset_status       : out std_logic;                                         --            hip_rst.reset_status
		serdes_pll_locked  : out std_logic;                                         --                   .serdes_pll_locked
		pld_clk_inuse      : out std_logic;                                         --                   .pld_clk_inuse
		pld_core_ready     : in  std_logic                      := '0';             --                   .pld_core_ready
		testin_zero        : out std_logic;                                         --                   .testin_zero
		reconfig_to_xcvr   : in  std_logic_vector(699 downto 0) := (others => '0'); --   reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr : out std_logic_vector(459 downto 0);                    -- reconfig_from_xcvr.reconfig_from_xcvr
		rx_in0             : in  std_logic                      := '0';             --         hip_serial.rx_in0
		rx_in1             : in  std_logic                      := '0';             --                   .rx_in1
		rx_in2             : in  std_logic                      := '0';             --                   .rx_in2
		rx_in3             : in  std_logic                      := '0';             --                   .rx_in3
		rx_in4             : in  std_logic                      := '0';             --                   .rx_in4
		rx_in5             : in  std_logic                      := '0';             --                   .rx_in5
		rx_in6             : in  std_logic                      := '0';             --                   .rx_in6
		rx_in7             : in  std_logic                      := '0';             --                   .rx_in7
		tx_out0            : out std_logic;                                         --                   .tx_out0
		tx_out1            : out std_logic;                                         --                   .tx_out1
		tx_out2            : out std_logic;                                         --                   .tx_out2
		tx_out3            : out std_logic;                                         --                   .tx_out3
		tx_out4            : out std_logic;                                         --                   .tx_out4
		tx_out5            : out std_logic;                                         --                   .tx_out5
		tx_out6            : out std_logic;                                         --                   .tx_out6
		tx_out7            : out std_logic;                                         --                   .tx_out7
		sim_pipe_pclk_in   : in  std_logic                      := '0';             --           hip_pipe.sim_pipe_pclk_in
		sim_pipe_rate      : out std_logic_vector(1 downto 0);                      --                   .sim_pipe_rate
		sim_ltssmstate     : out std_logic_vector(4 downto 0);                      --                   .sim_ltssmstate
		eidleinfersel0     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel0
		eidleinfersel1     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel1
		eidleinfersel2     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel2
		eidleinfersel3     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel3
		eidleinfersel4     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel4
		eidleinfersel5     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel5
		eidleinfersel6     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel6
		eidleinfersel7     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel7
		powerdown0         : out std_logic_vector(1 downto 0);                      --                   .powerdown0
		powerdown1         : out std_logic_vector(1 downto 0);                      --                   .powerdown1
		powerdown2         : out std_logic_vector(1 downto 0);                      --                   .powerdown2
		powerdown3         : out std_logic_vector(1 downto 0);                      --                   .powerdown3
		powerdown4         : out std_logic_vector(1 downto 0);                      --                   .powerdown4
		powerdown5         : out std_logic_vector(1 downto 0);                      --                   .powerdown5
		powerdown6         : out std_logic_vector(1 downto 0);                      --                   .powerdown6
		powerdown7         : out std_logic_vector(1 downto 0);                      --                   .powerdown7
		rxpolarity0        : out std_logic;                                         --                   .rxpolarity0
		rxpolarity1        : out std_logic;                                         --                   .rxpolarity1
		rxpolarity2        : out std_logic;                                         --                   .rxpolarity2
		rxpolarity3        : out std_logic;                                         --                   .rxpolarity3
		rxpolarity4        : out std_logic;                                         --                   .rxpolarity4
		rxpolarity5        : out std_logic;                                         --                   .rxpolarity5
		rxpolarity6        : out std_logic;                                         --                   .rxpolarity6
		rxpolarity7        : out std_logic;                                         --                   .rxpolarity7
		txcompl0           : out std_logic;                                         --                   .txcompl0
		txcompl1           : out std_logic;                                         --                   .txcompl1
		txcompl2           : out std_logic;                                         --                   .txcompl2
		txcompl3           : out std_logic;                                         --                   .txcompl3
		txcompl4           : out std_logic;                                         --                   .txcompl4
		txcompl5           : out std_logic;                                         --                   .txcompl5
		txcompl6           : out std_logic;                                         --                   .txcompl6
		txcompl7           : out std_logic;                                         --                   .txcompl7
		txdata0            : out std_logic_vector(7 downto 0);                      --                   .txdata0
		txdata1            : out std_logic_vector(7 downto 0);                      --                   .txdata1
		txdata2            : out std_logic_vector(7 downto 0);                      --                   .txdata2
		txdata3            : out std_logic_vector(7 downto 0);                      --                   .txdata3
		txdata4            : out std_logic_vector(7 downto 0);                      --                   .txdata4
		txdata5            : out std_logic_vector(7 downto 0);                      --                   .txdata5
		txdata6            : out std_logic_vector(7 downto 0);                      --                   .txdata6
		txdata7            : out std_logic_vector(7 downto 0);                      --                   .txdata7
		txdatak0           : out std_logic;                                         --                   .txdatak0
		txdatak1           : out std_logic;                                         --                   .txdatak1
		txdatak2           : out std_logic;                                         --                   .txdatak2
		txdatak3           : out std_logic;                                         --                   .txdatak3
		txdatak4           : out std_logic;                                         --                   .txdatak4
		txdatak5           : out std_logic;                                         --                   .txdatak5
		txdatak6           : out std_logic;                                         --                   .txdatak6
		txdatak7           : out std_logic;                                         --                   .txdatak7
		txdetectrx0        : out std_logic;                                         --                   .txdetectrx0
		txdetectrx1        : out std_logic;                                         --                   .txdetectrx1
		txdetectrx2        : out std_logic;                                         --                   .txdetectrx2
		txdetectrx3        : out std_logic;                                         --                   .txdetectrx3
		txdetectrx4        : out std_logic;                                         --                   .txdetectrx4
		txdetectrx5        : out std_logic;                                         --                   .txdetectrx5
		txdetectrx6        : out std_logic;                                         --                   .txdetectrx6
		txdetectrx7        : out std_logic;                                         --                   .txdetectrx7
		txelecidle0        : out std_logic;                                         --                   .txelecidle0
		txelecidle1        : out std_logic;                                         --                   .txelecidle1
		txelecidle2        : out std_logic;                                         --                   .txelecidle2
		txelecidle3        : out std_logic;                                         --                   .txelecidle3
		txelecidle4        : out std_logic;                                         --                   .txelecidle4
		txelecidle5        : out std_logic;                                         --                   .txelecidle5
		txelecidle6        : out std_logic;                                         --                   .txelecidle6
		txelecidle7        : out std_logic;                                         --                   .txelecidle7
		txdeemph0          : out std_logic;                                         --                   .txdeemph0
		txdeemph1          : out std_logic;                                         --                   .txdeemph1
		txdeemph2          : out std_logic;                                         --                   .txdeemph2
		txdeemph3          : out std_logic;                                         --                   .txdeemph3
		txdeemph4          : out std_logic;                                         --                   .txdeemph4
		txdeemph5          : out std_logic;                                         --                   .txdeemph5
		txdeemph6          : out std_logic;                                         --                   .txdeemph6
		txdeemph7          : out std_logic;                                         --                   .txdeemph7
		txmargin0          : out std_logic_vector(2 downto 0);                      --                   .txmargin0
		txmargin1          : out std_logic_vector(2 downto 0);                      --                   .txmargin1
		txmargin2          : out std_logic_vector(2 downto 0);                      --                   .txmargin2
		txmargin3          : out std_logic_vector(2 downto 0);                      --                   .txmargin3
		txmargin4          : out std_logic_vector(2 downto 0);                      --                   .txmargin4
		txmargin5          : out std_logic_vector(2 downto 0);                      --                   .txmargin5
		txmargin6          : out std_logic_vector(2 downto 0);                      --                   .txmargin6
		txmargin7          : out std_logic_vector(2 downto 0);                      --                   .txmargin7
		txswing0           : out std_logic;                                         --                   .txswing0
		txswing1           : out std_logic;                                         --                   .txswing1
		txswing2           : out std_logic;                                         --                   .txswing2
		txswing3           : out std_logic;                                         --                   .txswing3
		txswing4           : out std_logic;                                         --                   .txswing4
		txswing5           : out std_logic;                                         --                   .txswing5
		txswing6           : out std_logic;                                         --                   .txswing6
		txswing7           : out std_logic;                                         --                   .txswing7
		phystatus0         : in  std_logic                      := '0';             --                   .phystatus0
		phystatus1         : in  std_logic                      := '0';             --                   .phystatus1
		phystatus2         : in  std_logic                      := '0';             --                   .phystatus2
		phystatus3         : in  std_logic                      := '0';             --                   .phystatus3
		phystatus4         : in  std_logic                      := '0';             --                   .phystatus4
		phystatus5         : in  std_logic                      := '0';             --                   .phystatus5
		phystatus6         : in  std_logic                      := '0';             --                   .phystatus6
		phystatus7         : in  std_logic                      := '0';             --                   .phystatus7
		rxdata0            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata0
		rxdata1            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata1
		rxdata2            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata2
		rxdata3            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata3
		rxdata4            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata4
		rxdata5            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata5
		rxdata6            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata6
		rxdata7            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata7
		rxdatak0           : in  std_logic                      := '0';             --                   .rxdatak0
		rxdatak1           : in  std_logic                      := '0';             --                   .rxdatak1
		rxdatak2           : in  std_logic                      := '0';             --                   .rxdatak2
		rxdatak3           : in  std_logic                      := '0';             --                   .rxdatak3
		rxdatak4           : in  std_logic                      := '0';             --                   .rxdatak4
		rxdatak5           : in  std_logic                      := '0';             --                   .rxdatak5
		rxdatak6           : in  std_logic                      := '0';             --                   .rxdatak6
		rxdatak7           : in  std_logic                      := '0';             --                   .rxdatak7
		rxelecidle0        : in  std_logic                      := '0';             --                   .rxelecidle0
		rxelecidle1        : in  std_logic                      := '0';             --                   .rxelecidle1
		rxelecidle2        : in  std_logic                      := '0';             --                   .rxelecidle2
		rxelecidle3        : in  std_logic                      := '0';             --                   .rxelecidle3
		rxelecidle4        : in  std_logic                      := '0';             --                   .rxelecidle4
		rxelecidle5        : in  std_logic                      := '0';             --                   .rxelecidle5
		rxelecidle6        : in  std_logic                      := '0';             --                   .rxelecidle6
		rxelecidle7        : in  std_logic                      := '0';             --                   .rxelecidle7
		rxstatus0          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus0
		rxstatus1          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus1
		rxstatus2          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus2
		rxstatus3          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus3
		rxstatus4          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus4
		rxstatus5          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus5
		rxstatus6          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus6
		rxstatus7          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus7
		rxvalid0           : in  std_logic                      := '0';             --                   .rxvalid0
		rxvalid1           : in  std_logic                      := '0';             --                   .rxvalid1
		rxvalid2           : in  std_logic                      := '0';             --                   .rxvalid2
		rxvalid3           : in  std_logic                      := '0';             --                   .rxvalid3
		rxvalid4           : in  std_logic                      := '0';             --                   .rxvalid4
		rxvalid5           : in  std_logic                      := '0';             --                   .rxvalid5
		rxvalid6           : in  std_logic                      := '0';             --                   .rxvalid6
		rxvalid7           : in  std_logic                      := '0';             --                   .rxvalid7
		app_int_sts        : in  std_logic                      := '0';             --            int_msi.app_int_sts
		app_msi_num        : in  std_logic_vector(4 downto 0)   := (others => '0'); --                   .app_msi_num
		app_msi_req        : in  std_logic                      := '0';             --                   .app_msi_req
		app_msi_tc         : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .app_msi_tc
		app_int_ack        : out std_logic;                                         --                   .app_int_ack
		app_msi_ack        : out std_logic;                                         --                   .app_msi_ack
		test_in            : in  std_logic_vector(31 downto 0)  := (others => '0'); --           hip_ctrl.test_in
		simu_mode_pipe     : in  std_logic                      := '0';             --                   .simu_mode_pipe
		derr_cor_ext_rcv   : out std_logic;                                         --         hip_status.derr_cor_ext_rcv
		derr_cor_ext_rpl   : out std_logic;                                         --                   .derr_cor_ext_rpl
		derr_rpl           : out std_logic;                                         --                   .derr_rpl
		dlup               : out std_logic;                                         --                   .dlup
		dlup_exit          : out std_logic;                                         --                   .dlup_exit
		ev128ns            : out std_logic;                                         --                   .ev128ns
		ev1us              : out std_logic;                                         --                   .ev1us
		hotrst_exit        : out std_logic;                                         --                   .hotrst_exit
		int_status         : out std_logic_vector(3 downto 0);                      --                   .int_status
		l2_exit            : out std_logic;                                         --                   .l2_exit
		lane_act           : out std_logic_vector(3 downto 0);                      --                   .lane_act
		ltssmstate         : out std_logic_vector(4 downto 0);                      --                   .ltssmstate
		rx_par_err         : out std_logic;                                         --                   .rx_par_err
		tx_par_err         : out std_logic_vector(1 downto 0);                      --                   .tx_par_err
		cfg_par_err        : out std_logic;                                         --                   .cfg_par_err
		ko_cpl_spc_header  : out std_logic_vector(7 downto 0);                      --                   .ko_cpl_spc_header
		ko_cpl_spc_data    : out std_logic_vector(11 downto 0);                     --                   .ko_cpl_spc_data
		currentspeed       : out std_logic_vector(1 downto 0)                       --   hip_currentspeed.currentspeed
	);
end entity pcie_SV_hard_ip;

architecture rtl of pcie_SV_hard_ip is
	component altpcie_sv_hip_ast_hwtcl is
		generic (
			lane_mask_hwtcl                          : string  := "x4";
			gen123_lane_rate_mode_hwtcl              : string  := "Gen1 (2.5 Gbps)";
			port_type_hwtcl                          : string  := "Native endpoint";
			pcie_spec_version_hwtcl                  : string  := "2.1";
			ast_width_hwtcl                          : string  := "Avalon-ST 64-bit";
			pll_refclk_freq_hwtcl                    : string  := "100 MHz";
			set_pld_clk_x1_625MHz_hwtcl              : integer := 0;
			use_ast_parity                           : integer := 0;
			multiple_packets_per_cycle_hwtcl         : integer := 0;
			in_cvp_mode_hwtcl                        : integer := 0;
			use_pci_ext_hwtcl                        : integer := 0;
			use_pcie_ext_hwtcl                       : integer := 0;
			use_config_bypass_hwtcl                  : integer := 0;
			hip_reconfig_hwtcl                       : integer := 0;
			enable_tl_only_sim_hwtcl                 : integer := 0;
			bar0_size_mask_hwtcl                     : integer := 28;
			bar0_io_space_hwtcl                      : string  := "Disabled";
			bar0_64bit_mem_space_hwtcl               : string  := "Enabled";
			bar0_prefetchable_hwtcl                  : string  := "Enabled";
			bar1_size_mask_hwtcl                     : integer := 0;
			bar1_io_space_hwtcl                      : string  := "Disabled";
			bar1_prefetchable_hwtcl                  : string  := "Disabled";
			bar2_size_mask_hwtcl                     : integer := 0;
			bar2_io_space_hwtcl                      : string  := "Disabled";
			bar2_64bit_mem_space_hwtcl               : string  := "Disabled";
			bar2_prefetchable_hwtcl                  : string  := "Disabled";
			bar3_size_mask_hwtcl                     : integer := 0;
			bar3_io_space_hwtcl                      : string  := "Disabled";
			bar3_prefetchable_hwtcl                  : string  := "Disabled";
			bar4_size_mask_hwtcl                     : integer := 0;
			bar4_io_space_hwtcl                      : string  := "Disabled";
			bar4_64bit_mem_space_hwtcl               : string  := "Disabled";
			bar4_prefetchable_hwtcl                  : string  := "Disabled";
			bar5_size_mask_hwtcl                     : integer := 0;
			bar5_io_space_hwtcl                      : string  := "Disabled";
			bar5_prefetchable_hwtcl                  : string  := "Disabled";
			expansion_base_address_register_hwtcl    : integer := 0;
			io_window_addr_width_hwtcl               : integer := 0;
			prefetchable_mem_window_addr_width_hwtcl : integer := 0;
			vendor_id_hwtcl                          : integer := 0;
			device_id_hwtcl                          : integer := 1;
			revision_id_hwtcl                        : integer := 1;
			class_code_hwtcl                         : integer := 0;
			subsystem_vendor_id_hwtcl                : integer := 0;
			subsystem_device_id_hwtcl                : integer := 0;
			max_payload_size_hwtcl                   : integer := 128;
			extend_tag_field_hwtcl                   : string  := "32";
			completion_timeout_hwtcl                 : string  := "ABCD";
			enable_completion_timeout_disable_hwtcl  : integer := 1;
			use_aer_hwtcl                            : integer := 0;
			ecrc_check_capable_hwtcl                 : integer := 0;
			ecrc_gen_capable_hwtcl                   : integer := 0;
			use_crc_forwarding_hwtcl                 : integer := 0;
			port_link_number_hwtcl                   : integer := 1;
			dll_active_report_support_hwtcl          : integer := 0;
			surprise_down_error_support_hwtcl        : integer := 0;
			slotclkcfg_hwtcl                         : integer := 1;
			msi_multi_message_capable_hwtcl          : string  := "4";
			msi_64bit_addressing_capable_hwtcl       : string  := "true";
			msi_masking_capable_hwtcl                : string  := "false";
			msi_support_hwtcl                        : string  := "true";
			enable_function_msix_support_hwtcl       : integer := 0;
			msix_table_size_hwtcl                    : integer := 0;
			msix_table_offset_hwtcl                  : string  := "0";
			msix_table_bir_hwtcl                     : integer := 0;
			msix_pba_offset_hwtcl                    : string  := "0";
			msix_pba_bir_hwtcl                       : integer := 0;
			enable_slot_register_hwtcl               : integer := 0;
			slot_power_scale_hwtcl                   : integer := 0;
			slot_power_limit_hwtcl                   : integer := 0;
			slot_number_hwtcl                        : integer := 0;
			endpoint_l0_latency_hwtcl                : integer := 0;
			endpoint_l1_latency_hwtcl                : integer := 0;
			vsec_id_hwtcl                            : integer := 40960;
			vsec_rev_hwtcl                           : integer := 0;
			millisecond_cycle_count_hwtcl            : integer := 124250;
			port_width_be_hwtcl                      : integer := 8;
			port_width_data_hwtcl                    : integer := 64;
			gen3_dcbal_en_hwtcl                      : integer := 1;
			enable_pipe32_sim_hwtcl                  : integer := 0;
			fixed_preset_on                          : integer := 0;
			bypass_cdc_hwtcl                         : string  := "false";
			enable_rx_buffer_checking_hwtcl          : string  := "false";
			disable_link_x2_support_hwtcl            : string  := "false";
			wrong_device_id_hwtcl                    : string  := "disable";
			data_pack_rx_hwtcl                       : string  := "disable";
			ltssm_1ms_timeout_hwtcl                  : string  := "disable";
			ltssm_freqlocked_check_hwtcl             : string  := "disable";
			deskew_comma_hwtcl                       : string  := "skp_eieos_deskw";
			device_number_hwtcl                      : integer := 0;
			pipex1_debug_sel_hwtcl                   : string  := "disable";
			pclk_out_sel_hwtcl                       : string  := "pclk";
			no_soft_reset_hwtcl                      : string  := "false";
			maximum_current_hwtcl                    : integer := 0;
			d1_support_hwtcl                         : string  := "false";
			d2_support_hwtcl                         : string  := "false";
			d0_pme_hwtcl                             : string  := "false";
			d1_pme_hwtcl                             : string  := "false";
			d2_pme_hwtcl                             : string  := "false";
			d3_hot_pme_hwtcl                         : string  := "false";
			d3_cold_pme_hwtcl                        : string  := "false";
			low_priority_vc_hwtcl                    : string  := "single_vc";
			disable_snoop_packet_hwtcl               : string  := "false";
			enable_l1_aspm_hwtcl                     : string  := "false";
			rx_ei_l0s_hwtcl                          : integer := 0;
			enable_l0s_aspm_hwtcl                    : string  := "false";
			aspm_config_management_hwtcl             : string  := "false";
			l1_exit_latency_sameclock_hwtcl          : integer := 0;
			l1_exit_latency_diffclock_hwtcl          : integer := 0;
			hot_plug_support_hwtcl                   : integer := 0;
			extended_tag_reset_hwtcl                 : string  := "false";
			no_command_completed_hwtcl               : string  := "false";
			interrupt_pin_hwtcl                      : string  := "inta";
			bridge_port_vga_enable_hwtcl             : string  := "false";
			bridge_port_ssid_support_hwtcl           : string  := "false";
			ssvid_hwtcl                              : integer := 0;
			ssid_hwtcl                               : integer := 0;
			eie_before_nfts_count_hwtcl              : integer := 4;
			gen2_diffclock_nfts_count_hwtcl          : integer := 255;
			gen2_sameclock_nfts_count_hwtcl          : integer := 255;
			l0_exit_latency_sameclock_hwtcl          : integer := 6;
			l0_exit_latency_diffclock_hwtcl          : integer := 6;
			atomic_op_routing_hwtcl                  : string  := "false";
			atomic_op_completer_32bit_hwtcl          : string  := "false";
			atomic_op_completer_64bit_hwtcl          : string  := "false";
			cas_completer_128bit_hwtcl               : string  := "false";
			ltr_mechanism_hwtcl                      : string  := "false";
			tph_completer_hwtcl                      : string  := "false";
			extended_format_field_hwtcl              : string  := "false";
			atomic_malformed_hwtcl                   : string  := "true";
			flr_capability_hwtcl                     : string  := "false";
			enable_adapter_half_rate_mode_hwtcl      : string  := "false";
			vc0_clk_enable_hwtcl                     : string  := "true";
			register_pipe_signals_hwtcl              : string  := "false";
			skp_os_gen3_count_hwtcl                  : integer := 0;
			tx_cdc_almost_empty_hwtcl                : integer := 5;
			rx_l0s_count_idl_hwtcl                   : integer := 0;
			cdc_dummy_insert_limit_hwtcl             : integer := 11;
			ei_delay_powerdown_count_hwtcl           : integer := 10;
			skp_os_schedule_count_hwtcl              : integer := 0;
			fc_init_timer_hwtcl                      : integer := 1024;
			l01_entry_latency_hwtcl                  : integer := 31;
			flow_control_update_count_hwtcl          : integer := 30;
			flow_control_timeout_count_hwtcl         : integer := 200;
			retry_buffer_last_active_address_hwtcl   : integer := 2047;
			reserved_debug_hwtcl                     : integer := 0;
			bypass_clk_switch_hwtcl                  : string  := "true";
			l2_async_logic_hwtcl                     : string  := "disable";
			indicator_hwtcl                          : integer := 0;
			diffclock_nfts_count_hwtcl               : integer := 128;
			sameclock_nfts_count_hwtcl               : integer := 128;
			rx_cdc_almost_full_hwtcl                 : integer := 12;
			tx_cdc_almost_full_hwtcl                 : integer := 11;
			credit_buffer_allocation_aux_hwtcl       : string  := "balanced";
			vc0_rx_flow_ctrl_posted_header_hwtcl     : integer := 50;
			vc0_rx_flow_ctrl_posted_data_hwtcl       : integer := 358;
			vc0_rx_flow_ctrl_nonposted_header_hwtcl  : integer := 56;
			vc0_rx_flow_ctrl_nonposted_data_hwtcl    : integer := 0;
			vc0_rx_flow_ctrl_compl_header_hwtcl      : integer := 0;
			vc0_rx_flow_ctrl_compl_data_hwtcl        : integer := 0;
			cpl_spc_header_hwtcl                     : integer := 112;
			cpl_spc_data_hwtcl                       : integer := 448;
			gen3_rxfreqlock_counter_hwtcl            : integer := 0;
			gen3_skip_ph2_ph3_hwtcl                  : integer := 0;
			g3_bypass_equlz_hwtcl                    : integer := 0;
			cvp_data_compressed_hwtcl                : string  := "false";
			cvp_data_encrypted_hwtcl                 : string  := "false";
			cvp_mode_reset_hwtcl                     : string  := "false";
			cvp_clk_reset_hwtcl                      : string  := "false";
			cseb_cpl_status_during_cvp_hwtcl         : string  := "config_retry_status";
			core_clk_sel_hwtcl                       : string  := "pld_clk";
			cvp_rate_sel_hwtcl                       : string  := "full_rate";
			g3_dis_rx_use_prst_hwtcl                 : string  := "true";
			g3_dis_rx_use_prst_ep_hwtcl              : string  := "true";
			deemphasis_enable_hwtcl                  : string  := "false";
			reconfig_to_xcvr_width                   : integer := 10;
			reconfig_from_xcvr_width                 : integer := 10;
			single_rx_detect_hwtcl                   : integer := 0;
			hip_hard_reset_hwtcl                     : integer := 1;
			hwtcl_override_g2_txvod                  : integer := 1;
			rpre_emph_a_val_hwtcl                    : integer := 9;
			rpre_emph_b_val_hwtcl                    : integer := 0;
			rpre_emph_c_val_hwtcl                    : integer := 16;
			rpre_emph_d_val_hwtcl                    : integer := 13;
			rpre_emph_e_val_hwtcl                    : integer := 5;
			rvod_sel_a_val_hwtcl                     : integer := 42;
			rvod_sel_b_val_hwtcl                     : integer := 38;
			rvod_sel_c_val_hwtcl                     : integer := 38;
			rvod_sel_d_val_hwtcl                     : integer := 43;
			rvod_sel_e_val_hwtcl                     : integer := 15;
			hwtcl_override_g3rxcoef                  : integer := 0;
			gen3_coeff_1_hwtcl                       : integer := 7;
			gen3_coeff_1_sel_hwtcl                   : string  := "preset_1";
			gen3_coeff_1_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_1_nxtber_more_ptr_hwtcl       : integer := 1;
			gen3_coeff_1_nxtber_more_hwtcl           : string  := "g3_coeff_1_nxtber_more";
			gen3_coeff_1_nxtber_less_ptr_hwtcl       : integer := 1;
			gen3_coeff_1_nxtber_less_hwtcl           : string  := "g3_coeff_1_nxtber_less";
			gen3_coeff_1_reqber_hwtcl                : integer := 0;
			gen3_coeff_1_ber_meas_hwtcl              : integer := 2;
			gen3_coeff_2_hwtcl                       : integer := 0;
			gen3_coeff_2_sel_hwtcl                   : string  := "preset_2";
			gen3_coeff_2_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_2_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_2_nxtber_more_hwtcl           : string  := "g3_coeff_2_nxtber_more";
			gen3_coeff_2_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_2_nxtber_less_hwtcl           : string  := "g3_coeff_2_nxtber_less";
			gen3_coeff_2_reqber_hwtcl                : integer := 0;
			gen3_coeff_2_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_3_hwtcl                       : integer := 0;
			gen3_coeff_3_sel_hwtcl                   : string  := "preset_3";
			gen3_coeff_3_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_3_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_3_nxtber_more_hwtcl           : string  := "g3_coeff_3_nxtber_more";
			gen3_coeff_3_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_3_nxtber_less_hwtcl           : string  := "g3_coeff_3_nxtber_less";
			gen3_coeff_3_reqber_hwtcl                : integer := 0;
			gen3_coeff_3_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_4_hwtcl                       : integer := 0;
			gen3_coeff_4_sel_hwtcl                   : string  := "preset_4";
			gen3_coeff_4_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_4_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_4_nxtber_more_hwtcl           : string  := "g3_coeff_4_nxtber_more";
			gen3_coeff_4_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_4_nxtber_less_hwtcl           : string  := "g3_coeff_4_nxtber_less";
			gen3_coeff_4_reqber_hwtcl                : integer := 0;
			gen3_coeff_4_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_5_hwtcl                       : integer := 0;
			gen3_coeff_5_sel_hwtcl                   : string  := "preset_5";
			gen3_coeff_5_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_5_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_5_nxtber_more_hwtcl           : string  := "g3_coeff_5_nxtber_more";
			gen3_coeff_5_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_5_nxtber_less_hwtcl           : string  := "g3_coeff_5_nxtber_less";
			gen3_coeff_5_reqber_hwtcl                : integer := 0;
			gen3_coeff_5_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_6_hwtcl                       : integer := 0;
			gen3_coeff_6_sel_hwtcl                   : string  := "preset_6";
			gen3_coeff_6_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_6_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_6_nxtber_more_hwtcl           : string  := "g3_coeff_6_nxtber_more";
			gen3_coeff_6_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_6_nxtber_less_hwtcl           : string  := "g3_coeff_6_nxtber_less";
			gen3_coeff_6_reqber_hwtcl                : integer := 0;
			gen3_coeff_6_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_7_hwtcl                       : integer := 0;
			gen3_coeff_7_sel_hwtcl                   : string  := "preset_7";
			gen3_coeff_7_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_7_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_7_nxtber_more_hwtcl           : string  := "g3_coeff_7_nxtber_more";
			gen3_coeff_7_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_7_nxtber_less_hwtcl           : string  := "g3_coeff_7_nxtber_less";
			gen3_coeff_7_reqber_hwtcl                : integer := 0;
			gen3_coeff_7_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_8_hwtcl                       : integer := 0;
			gen3_coeff_8_sel_hwtcl                   : string  := "preset_8";
			gen3_coeff_8_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_8_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_8_nxtber_more_hwtcl           : string  := "g3_coeff_8_nxtber_more";
			gen3_coeff_8_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_8_nxtber_less_hwtcl           : string  := "g3_coeff_8_nxtber_less";
			gen3_coeff_8_reqber_hwtcl                : integer := 0;
			gen3_coeff_8_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_9_hwtcl                       : integer := 0;
			gen3_coeff_9_sel_hwtcl                   : string  := "preset_9";
			gen3_coeff_9_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_9_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_9_nxtber_more_hwtcl           : string  := "g3_coeff_9_nxtber_more";
			gen3_coeff_9_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_9_nxtber_less_hwtcl           : string  := "g3_coeff_9_nxtber_less";
			gen3_coeff_9_reqber_hwtcl                : integer := 0;
			gen3_coeff_9_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_10_hwtcl                      : integer := 0;
			gen3_coeff_10_sel_hwtcl                  : string  := "preset_10";
			gen3_coeff_10_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_10_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_10_nxtber_more_hwtcl          : string  := "g3_coeff_10_nxtber_more";
			gen3_coeff_10_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_10_nxtber_less_hwtcl          : string  := "g3_coeff_10_nxtber_less";
			gen3_coeff_10_reqber_hwtcl               : integer := 0;
			gen3_coeff_10_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_11_hwtcl                      : integer := 0;
			gen3_coeff_11_sel_hwtcl                  : string  := "preset_11";
			gen3_coeff_11_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_11_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_11_nxtber_more_hwtcl          : string  := "g3_coeff_11_nxtber_more";
			gen3_coeff_11_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_11_nxtber_less_hwtcl          : string  := "g3_coeff_11_nxtber_less";
			gen3_coeff_11_reqber_hwtcl               : integer := 0;
			gen3_coeff_11_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_12_hwtcl                      : integer := 0;
			gen3_coeff_12_sel_hwtcl                  : string  := "preset_12";
			gen3_coeff_12_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_12_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_12_nxtber_more_hwtcl          : string  := "g3_coeff_12_nxtber_more";
			gen3_coeff_12_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_12_nxtber_less_hwtcl          : string  := "g3_coeff_12_nxtber_less";
			gen3_coeff_12_reqber_hwtcl               : integer := 0;
			gen3_coeff_12_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_13_hwtcl                      : integer := 0;
			gen3_coeff_13_sel_hwtcl                  : string  := "preset_13";
			gen3_coeff_13_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_13_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_13_nxtber_more_hwtcl          : string  := "g3_coeff_13_nxtber_more";
			gen3_coeff_13_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_13_nxtber_less_hwtcl          : string  := "g3_coeff_13_nxtber_less";
			gen3_coeff_13_reqber_hwtcl               : integer := 0;
			gen3_coeff_13_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_14_hwtcl                      : integer := 0;
			gen3_coeff_14_sel_hwtcl                  : string  := "preset_14";
			gen3_coeff_14_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_14_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_14_nxtber_more_hwtcl          : string  := "g3_coeff_14_nxtber_more";
			gen3_coeff_14_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_14_nxtber_less_hwtcl          : string  := "g3_coeff_14_nxtber_less";
			gen3_coeff_14_reqber_hwtcl               : integer := 0;
			gen3_coeff_14_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_15_hwtcl                      : integer := 0;
			gen3_coeff_15_sel_hwtcl                  : string  := "preset_15";
			gen3_coeff_15_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_15_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_15_nxtber_more_hwtcl          : string  := "g3_coeff_15_nxtber_more";
			gen3_coeff_15_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_15_nxtber_less_hwtcl          : string  := "g3_coeff_15_nxtber_less";
			gen3_coeff_15_reqber_hwtcl               : integer := 0;
			gen3_coeff_15_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_16_hwtcl                      : integer := 0;
			gen3_coeff_16_sel_hwtcl                  : string  := "preset_16";
			gen3_coeff_16_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_16_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_16_nxtber_more_hwtcl          : string  := "g3_coeff_16_nxtber_more";
			gen3_coeff_16_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_16_nxtber_less_hwtcl          : string  := "g3_coeff_16_nxtber_less";
			gen3_coeff_16_reqber_hwtcl               : integer := 0;
			gen3_coeff_16_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_17_hwtcl                      : integer := 0;
			gen3_coeff_17_sel_hwtcl                  : string  := "preset_17";
			gen3_coeff_17_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_17_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_17_nxtber_more_hwtcl          : string  := "g3_coeff_17_nxtber_more";
			gen3_coeff_17_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_17_nxtber_less_hwtcl          : string  := "g3_coeff_17_nxtber_less";
			gen3_coeff_17_reqber_hwtcl               : integer := 0;
			gen3_coeff_17_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_18_hwtcl                      : integer := 0;
			gen3_coeff_18_sel_hwtcl                  : string  := "preset_18";
			gen3_coeff_18_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_18_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_18_nxtber_more_hwtcl          : string  := "g3_coeff_18_nxtber_more";
			gen3_coeff_18_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_18_nxtber_less_hwtcl          : string  := "g3_coeff_18_nxtber_less";
			gen3_coeff_18_reqber_hwtcl               : integer := 0;
			gen3_coeff_18_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_19_hwtcl                      : integer := 0;
			gen3_coeff_19_sel_hwtcl                  : string  := "preset_19";
			gen3_coeff_19_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_19_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_19_nxtber_more_hwtcl          : string  := "g3_coeff_19_nxtber_more";
			gen3_coeff_19_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_19_nxtber_less_hwtcl          : string  := "g3_coeff_19_nxtber_less";
			gen3_coeff_19_reqber_hwtcl               : integer := 0;
			gen3_coeff_19_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_20_hwtcl                      : integer := 0;
			gen3_coeff_20_sel_hwtcl                  : string  := "preset_20";
			gen3_coeff_20_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_20_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_20_nxtber_more_hwtcl          : string  := "g3_coeff_20_nxtber_more";
			gen3_coeff_20_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_20_nxtber_less_hwtcl          : string  := "g3_coeff_20_nxtber_less";
			gen3_coeff_20_reqber_hwtcl               : integer := 0;
			gen3_coeff_20_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_21_hwtcl                      : integer := 0;
			gen3_coeff_21_sel_hwtcl                  : string  := "preset_21";
			gen3_coeff_21_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_21_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_21_nxtber_more_hwtcl          : string  := "g3_coeff_21_nxtber_more";
			gen3_coeff_21_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_21_nxtber_less_hwtcl          : string  := "g3_coeff_21_nxtber_less";
			gen3_coeff_21_reqber_hwtcl               : integer := 0;
			gen3_coeff_21_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_22_hwtcl                      : integer := 0;
			gen3_coeff_22_sel_hwtcl                  : string  := "preset_22";
			gen3_coeff_22_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_22_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_22_nxtber_more_hwtcl          : string  := "g3_coeff_22_nxtber_more";
			gen3_coeff_22_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_22_nxtber_less_hwtcl          : string  := "g3_coeff_22_nxtber_less";
			gen3_coeff_22_reqber_hwtcl               : integer := 0;
			gen3_coeff_22_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_23_hwtcl                      : integer := 0;
			gen3_coeff_23_sel_hwtcl                  : string  := "preset_23";
			gen3_coeff_23_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_23_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_23_nxtber_more_hwtcl          : string  := "g3_coeff_23_nxtber_more";
			gen3_coeff_23_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_23_nxtber_less_hwtcl          : string  := "g3_coeff_23_nxtber_less";
			gen3_coeff_23_reqber_hwtcl               : integer := 0;
			gen3_coeff_23_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_24_hwtcl                      : integer := 0;
			gen3_coeff_24_sel_hwtcl                  : string  := "preset_24";
			gen3_coeff_24_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_24_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_24_nxtber_more_hwtcl          : string  := "g3_coeff_24_nxtber_more";
			gen3_coeff_24_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_24_nxtber_less_hwtcl          : string  := "g3_coeff_24_nxtber_less";
			gen3_coeff_24_reqber_hwtcl               : integer := 0;
			gen3_coeff_24_ber_meas_hwtcl             : integer := 0;
			hwtcl_override_g3txcoef                  : integer := 0;
			gen3_preset_coeff_1_hwtcl                : integer := 0;
			gen3_preset_coeff_2_hwtcl                : integer := 0;
			gen3_preset_coeff_3_hwtcl                : integer := 0;
			gen3_preset_coeff_4_hwtcl                : integer := 0;
			gen3_preset_coeff_5_hwtcl                : integer := 0;
			gen3_preset_coeff_6_hwtcl                : integer := 0;
			gen3_preset_coeff_7_hwtcl                : integer := 0;
			gen3_preset_coeff_8_hwtcl                : integer := 0;
			gen3_preset_coeff_9_hwtcl                : integer := 0;
			gen3_preset_coeff_10_hwtcl               : integer := 0;
			gen3_preset_coeff_11_hwtcl               : integer := 0;
			gen3_low_freq_hwtcl                      : integer := 0;
			full_swing_hwtcl                         : integer := 35;
			gen3_full_swing_hwtcl                    : integer := 35;
			use_atx_pll_hwtcl                        : integer := 0;
			low_latency_mode_hwtcl                   : integer := 0
		);
		port (
			npor                   : in  std_logic                       := 'X';             -- npor
			pin_perst              : in  std_logic                       := 'X';             -- pin_perst
			lmi_addr               : in  std_logic_vector(11 downto 0)   := (others => 'X'); -- lmi_addr
			lmi_din                : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- lmi_din
			lmi_rden               : in  std_logic                       := 'X';             -- lmi_rden
			lmi_wren               : in  std_logic                       := 'X';             -- lmi_wren
			lmi_ack                : out std_logic;                                          -- lmi_ack
			lmi_dout               : out std_logic_vector(31 downto 0);                      -- lmi_dout
			hpg_ctrler             : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- hpg_ctrler
			tl_cfg_add             : out std_logic_vector(3 downto 0);                       -- tl_cfg_add
			tl_cfg_ctl             : out std_logic_vector(31 downto 0);                      -- tl_cfg_ctl
			tl_cfg_sts             : out std_logic_vector(52 downto 0);                      -- tl_cfg_sts
			cpl_err                : in  std_logic_vector(6 downto 0)    := (others => 'X'); -- cpl_err
			cpl_pending            : in  std_logic                       := 'X';             -- cpl_pending
			pm_auxpwr              : in  std_logic                       := 'X';             -- pm_auxpwr
			pm_data                : in  std_logic_vector(9 downto 0)    := (others => 'X'); -- pm_data
			pme_to_cr              : in  std_logic                       := 'X';             -- pme_to_cr
			pm_event               : in  std_logic                       := 'X';             -- pm_event
			pme_to_sr              : out std_logic;                                          -- pme_to_sr
			rx_st_sop              : out std_logic_vector(0 downto 0);                       -- startofpacket
			rx_st_eop              : out std_logic_vector(0 downto 0);                       -- endofpacket
			rx_st_err              : out std_logic_vector(0 downto 0);                       -- error
			rx_st_valid            : out std_logic_vector(0 downto 0);                       -- valid
			rx_st_empty            : out std_logic_vector(1 downto 0);                       -- empty
			rx_st_ready            : in  std_logic                       := 'X';             -- ready
			rx_st_data             : out std_logic_vector(127 downto 0);                     -- data
			rx_st_bar              : out std_logic_vector(7 downto 0);                       -- rx_st_bar
			rx_st_mask             : in  std_logic                       := 'X';             -- rx_st_mask
			tx_st_sop              : in  std_logic_vector(0 downto 0)    := (others => 'X'); -- startofpacket
			tx_st_eop              : in  std_logic_vector(0 downto 0)    := (others => 'X'); -- endofpacket
			tx_st_err              : in  std_logic_vector(0 downto 0)    := (others => 'X'); -- error
			tx_st_valid            : in  std_logic_vector(0 downto 0)    := (others => 'X'); -- valid
			tx_st_empty            : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- empty
			tx_st_ready            : out std_logic;                                          -- ready
			tx_st_data             : in  std_logic_vector(127 downto 0)  := (others => 'X'); -- data
			tx_cred_datafccp       : out std_logic_vector(11 downto 0);                      -- tx_cred_datafccp
			tx_cred_datafcnp       : out std_logic_vector(11 downto 0);                      -- tx_cred_datafcnp
			tx_cred_datafcp        : out std_logic_vector(11 downto 0);                      -- tx_cred_datafcp
			tx_cred_fchipcons      : out std_logic_vector(5 downto 0);                       -- tx_cred_fchipcons
			tx_cred_fcinfinite     : out std_logic_vector(5 downto 0);                       -- tx_cred_fcinfinite
			tx_cred_hdrfccp        : out std_logic_vector(7 downto 0);                       -- tx_cred_hdrfccp
			tx_cred_hdrfcnp        : out std_logic_vector(7 downto 0);                       -- tx_cred_hdrfcnp
			tx_cred_hdrfcp         : out std_logic_vector(7 downto 0);                       -- tx_cred_hdrfcp
			pld_clk                : in  std_logic                       := 'X';             -- clk
			coreclkout_hip         : out std_logic;                                          -- clk
			refclk                 : in  std_logic                       := 'X';             -- clk
			reset_status           : out std_logic;                                          -- reset_status
			serdes_pll_locked      : out std_logic;                                          -- serdes_pll_locked
			pld_clk_inuse          : out std_logic;                                          -- pld_clk_inuse
			pld_core_ready         : in  std_logic                       := 'X';             -- pld_core_ready
			testin_zero            : out std_logic;                                          -- testin_zero
			reconfig_to_xcvr       : in  std_logic_vector(699 downto 0)  := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr     : out std_logic_vector(459 downto 0);                     -- reconfig_from_xcvr
			rx_in0                 : in  std_logic                       := 'X';             -- rx_in0
			rx_in1                 : in  std_logic                       := 'X';             -- rx_in1
			rx_in2                 : in  std_logic                       := 'X';             -- rx_in2
			rx_in3                 : in  std_logic                       := 'X';             -- rx_in3
			rx_in4                 : in  std_logic                       := 'X';             -- rx_in4
			rx_in5                 : in  std_logic                       := 'X';             -- rx_in5
			rx_in6                 : in  std_logic                       := 'X';             -- rx_in6
			rx_in7                 : in  std_logic                       := 'X';             -- rx_in7
			tx_out0                : out std_logic;                                          -- tx_out0
			tx_out1                : out std_logic;                                          -- tx_out1
			tx_out2                : out std_logic;                                          -- tx_out2
			tx_out3                : out std_logic;                                          -- tx_out3
			tx_out4                : out std_logic;                                          -- tx_out4
			tx_out5                : out std_logic;                                          -- tx_out5
			tx_out6                : out std_logic;                                          -- tx_out6
			tx_out7                : out std_logic;                                          -- tx_out7
			sim_pipe_pclk_in       : in  std_logic                       := 'X';             -- sim_pipe_pclk_in
			sim_pipe_rate          : out std_logic_vector(1 downto 0);                       -- sim_pipe_rate
			sim_ltssmstate         : out std_logic_vector(4 downto 0);                       -- sim_ltssmstate
			eidleinfersel0         : out std_logic_vector(2 downto 0);                       -- eidleinfersel0
			eidleinfersel1         : out std_logic_vector(2 downto 0);                       -- eidleinfersel1
			eidleinfersel2         : out std_logic_vector(2 downto 0);                       -- eidleinfersel2
			eidleinfersel3         : out std_logic_vector(2 downto 0);                       -- eidleinfersel3
			eidleinfersel4         : out std_logic_vector(2 downto 0);                       -- eidleinfersel4
			eidleinfersel5         : out std_logic_vector(2 downto 0);                       -- eidleinfersel5
			eidleinfersel6         : out std_logic_vector(2 downto 0);                       -- eidleinfersel6
			eidleinfersel7         : out std_logic_vector(2 downto 0);                       -- eidleinfersel7
			powerdown0             : out std_logic_vector(1 downto 0);                       -- powerdown0
			powerdown1             : out std_logic_vector(1 downto 0);                       -- powerdown1
			powerdown2             : out std_logic_vector(1 downto 0);                       -- powerdown2
			powerdown3             : out std_logic_vector(1 downto 0);                       -- powerdown3
			powerdown4             : out std_logic_vector(1 downto 0);                       -- powerdown4
			powerdown5             : out std_logic_vector(1 downto 0);                       -- powerdown5
			powerdown6             : out std_logic_vector(1 downto 0);                       -- powerdown6
			powerdown7             : out std_logic_vector(1 downto 0);                       -- powerdown7
			rxpolarity0            : out std_logic;                                          -- rxpolarity0
			rxpolarity1            : out std_logic;                                          -- rxpolarity1
			rxpolarity2            : out std_logic;                                          -- rxpolarity2
			rxpolarity3            : out std_logic;                                          -- rxpolarity3
			rxpolarity4            : out std_logic;                                          -- rxpolarity4
			rxpolarity5            : out std_logic;                                          -- rxpolarity5
			rxpolarity6            : out std_logic;                                          -- rxpolarity6
			rxpolarity7            : out std_logic;                                          -- rxpolarity7
			txcompl0               : out std_logic;                                          -- txcompl0
			txcompl1               : out std_logic;                                          -- txcompl1
			txcompl2               : out std_logic;                                          -- txcompl2
			txcompl3               : out std_logic;                                          -- txcompl3
			txcompl4               : out std_logic;                                          -- txcompl4
			txcompl5               : out std_logic;                                          -- txcompl5
			txcompl6               : out std_logic;                                          -- txcompl6
			txcompl7               : out std_logic;                                          -- txcompl7
			txdata0                : out std_logic_vector(7 downto 0);                       -- txdata0
			txdata1                : out std_logic_vector(7 downto 0);                       -- txdata1
			txdata2                : out std_logic_vector(7 downto 0);                       -- txdata2
			txdata3                : out std_logic_vector(7 downto 0);                       -- txdata3
			txdata4                : out std_logic_vector(7 downto 0);                       -- txdata4
			txdata5                : out std_logic_vector(7 downto 0);                       -- txdata5
			txdata6                : out std_logic_vector(7 downto 0);                       -- txdata6
			txdata7                : out std_logic_vector(7 downto 0);                       -- txdata7
			txdatak0               : out std_logic;                                          -- txdatak0
			txdatak1               : out std_logic;                                          -- txdatak1
			txdatak2               : out std_logic;                                          -- txdatak2
			txdatak3               : out std_logic;                                          -- txdatak3
			txdatak4               : out std_logic;                                          -- txdatak4
			txdatak5               : out std_logic;                                          -- txdatak5
			txdatak6               : out std_logic;                                          -- txdatak6
			txdatak7               : out std_logic;                                          -- txdatak7
			txdetectrx0            : out std_logic;                                          -- txdetectrx0
			txdetectrx1            : out std_logic;                                          -- txdetectrx1
			txdetectrx2            : out std_logic;                                          -- txdetectrx2
			txdetectrx3            : out std_logic;                                          -- txdetectrx3
			txdetectrx4            : out std_logic;                                          -- txdetectrx4
			txdetectrx5            : out std_logic;                                          -- txdetectrx5
			txdetectrx6            : out std_logic;                                          -- txdetectrx6
			txdetectrx7            : out std_logic;                                          -- txdetectrx7
			txelecidle0            : out std_logic;                                          -- txelecidle0
			txelecidle1            : out std_logic;                                          -- txelecidle1
			txelecidle2            : out std_logic;                                          -- txelecidle2
			txelecidle3            : out std_logic;                                          -- txelecidle3
			txelecidle4            : out std_logic;                                          -- txelecidle4
			txelecidle5            : out std_logic;                                          -- txelecidle5
			txelecidle6            : out std_logic;                                          -- txelecidle6
			txelecidle7            : out std_logic;                                          -- txelecidle7
			txdeemph0              : out std_logic;                                          -- txdeemph0
			txdeemph1              : out std_logic;                                          -- txdeemph1
			txdeemph2              : out std_logic;                                          -- txdeemph2
			txdeemph3              : out std_logic;                                          -- txdeemph3
			txdeemph4              : out std_logic;                                          -- txdeemph4
			txdeemph5              : out std_logic;                                          -- txdeemph5
			txdeemph6              : out std_logic;                                          -- txdeemph6
			txdeemph7              : out std_logic;                                          -- txdeemph7
			txmargin0              : out std_logic_vector(2 downto 0);                       -- txmargin0
			txmargin1              : out std_logic_vector(2 downto 0);                       -- txmargin1
			txmargin2              : out std_logic_vector(2 downto 0);                       -- txmargin2
			txmargin3              : out std_logic_vector(2 downto 0);                       -- txmargin3
			txmargin4              : out std_logic_vector(2 downto 0);                       -- txmargin4
			txmargin5              : out std_logic_vector(2 downto 0);                       -- txmargin5
			txmargin6              : out std_logic_vector(2 downto 0);                       -- txmargin6
			txmargin7              : out std_logic_vector(2 downto 0);                       -- txmargin7
			txswing0               : out std_logic;                                          -- txswing0
			txswing1               : out std_logic;                                          -- txswing1
			txswing2               : out std_logic;                                          -- txswing2
			txswing3               : out std_logic;                                          -- txswing3
			txswing4               : out std_logic;                                          -- txswing4
			txswing5               : out std_logic;                                          -- txswing5
			txswing6               : out std_logic;                                          -- txswing6
			txswing7               : out std_logic;                                          -- txswing7
			phystatus0             : in  std_logic                       := 'X';             -- phystatus0
			phystatus1             : in  std_logic                       := 'X';             -- phystatus1
			phystatus2             : in  std_logic                       := 'X';             -- phystatus2
			phystatus3             : in  std_logic                       := 'X';             -- phystatus3
			phystatus4             : in  std_logic                       := 'X';             -- phystatus4
			phystatus5             : in  std_logic                       := 'X';             -- phystatus5
			phystatus6             : in  std_logic                       := 'X';             -- phystatus6
			phystatus7             : in  std_logic                       := 'X';             -- phystatus7
			rxdata0                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata0
			rxdata1                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata1
			rxdata2                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata2
			rxdata3                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata3
			rxdata4                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata4
			rxdata5                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata5
			rxdata6                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata6
			rxdata7                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata7
			rxdatak0               : in  std_logic                       := 'X';             -- rxdatak0
			rxdatak1               : in  std_logic                       := 'X';             -- rxdatak1
			rxdatak2               : in  std_logic                       := 'X';             -- rxdatak2
			rxdatak3               : in  std_logic                       := 'X';             -- rxdatak3
			rxdatak4               : in  std_logic                       := 'X';             -- rxdatak4
			rxdatak5               : in  std_logic                       := 'X';             -- rxdatak5
			rxdatak6               : in  std_logic                       := 'X';             -- rxdatak6
			rxdatak7               : in  std_logic                       := 'X';             -- rxdatak7
			rxelecidle0            : in  std_logic                       := 'X';             -- rxelecidle0
			rxelecidle1            : in  std_logic                       := 'X';             -- rxelecidle1
			rxelecidle2            : in  std_logic                       := 'X';             -- rxelecidle2
			rxelecidle3            : in  std_logic                       := 'X';             -- rxelecidle3
			rxelecidle4            : in  std_logic                       := 'X';             -- rxelecidle4
			rxelecidle5            : in  std_logic                       := 'X';             -- rxelecidle5
			rxelecidle6            : in  std_logic                       := 'X';             -- rxelecidle6
			rxelecidle7            : in  std_logic                       := 'X';             -- rxelecidle7
			rxstatus0              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus0
			rxstatus1              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus1
			rxstatus2              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus2
			rxstatus3              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus3
			rxstatus4              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus4
			rxstatus5              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus5
			rxstatus6              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus6
			rxstatus7              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus7
			rxvalid0               : in  std_logic                       := 'X';             -- rxvalid0
			rxvalid1               : in  std_logic                       := 'X';             -- rxvalid1
			rxvalid2               : in  std_logic                       := 'X';             -- rxvalid2
			rxvalid3               : in  std_logic                       := 'X';             -- rxvalid3
			rxvalid4               : in  std_logic                       := 'X';             -- rxvalid4
			rxvalid5               : in  std_logic                       := 'X';             -- rxvalid5
			rxvalid6               : in  std_logic                       := 'X';             -- rxvalid6
			rxvalid7               : in  std_logic                       := 'X';             -- rxvalid7
			app_int_sts            : in  std_logic                       := 'X';             -- app_int_sts
			app_msi_num            : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- app_msi_num
			app_msi_req            : in  std_logic                       := 'X';             -- app_msi_req
			app_msi_tc             : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- app_msi_tc
			app_int_ack            : out std_logic;                                          -- app_int_ack
			app_msi_ack            : out std_logic;                                          -- app_msi_ack
			test_in                : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- test_in
			simu_mode_pipe         : in  std_logic                       := 'X';             -- simu_mode_pipe
			derr_cor_ext_rcv       : out std_logic;                                          -- derr_cor_ext_rcv
			derr_cor_ext_rpl       : out std_logic;                                          -- derr_cor_ext_rpl
			derr_rpl               : out std_logic;                                          -- derr_rpl
			dlup                   : out std_logic;                                          -- dlup
			dlup_exit              : out std_logic;                                          -- dlup_exit
			ev128ns                : out std_logic;                                          -- ev128ns
			ev1us                  : out std_logic;                                          -- ev1us
			hotrst_exit            : out std_logic;                                          -- hotrst_exit
			int_status             : out std_logic_vector(3 downto 0);                       -- int_status
			l2_exit                : out std_logic;                                          -- l2_exit
			lane_act               : out std_logic_vector(3 downto 0);                       -- lane_act
			ltssmstate             : out std_logic_vector(4 downto 0);                       -- ltssmstate
			rx_par_err             : out std_logic;                                          -- rx_par_err
			tx_par_err             : out std_logic_vector(1 downto 0);                       -- tx_par_err
			cfg_par_err            : out std_logic;                                          -- cfg_par_err
			ko_cpl_spc_header      : out std_logic_vector(7 downto 0);                       -- ko_cpl_spc_header
			ko_cpl_spc_data        : out std_logic_vector(11 downto 0);                      -- ko_cpl_spc_data
			currentspeed           : out std_logic_vector(1 downto 0);                       -- currentspeed
			rx_st_parity           : out std_logic_vector(15 downto 0);                      -- rx_st_parity
			rx_st_be               : out std_logic_vector(15 downto 0);                      -- rx_st_be
			tx_st_parity           : in  std_logic_vector(15 downto 0)   := (others => 'X'); -- tx_st_parity
			tx_cons_cred_sel       : in  std_logic                       := 'X';             -- tx_cons_cred_sel
			sim_pipe_pclk_out      : out std_logic;                                          -- sim_pipe_pclk_out
			rxdataskip0            : in  std_logic                       := 'X';             -- rxdataskip0
			rxdataskip1            : in  std_logic                       := 'X';             -- rxdataskip1
			rxdataskip2            : in  std_logic                       := 'X';             -- rxdataskip2
			rxdataskip3            : in  std_logic                       := 'X';             -- rxdataskip3
			rxdataskip4            : in  std_logic                       := 'X';             -- rxdataskip4
			rxdataskip5            : in  std_logic                       := 'X';             -- rxdataskip5
			rxdataskip6            : in  std_logic                       := 'X';             -- rxdataskip6
			rxdataskip7            : in  std_logic                       := 'X';             -- rxdataskip7
			rxblkst0               : in  std_logic                       := 'X';             -- rxblkst0
			rxblkst1               : in  std_logic                       := 'X';             -- rxblkst1
			rxblkst2               : in  std_logic                       := 'X';             -- rxblkst2
			rxblkst3               : in  std_logic                       := 'X';             -- rxblkst3
			rxblkst4               : in  std_logic                       := 'X';             -- rxblkst4
			rxblkst5               : in  std_logic                       := 'X';             -- rxblkst5
			rxblkst6               : in  std_logic                       := 'X';             -- rxblkst6
			rxblkst7               : in  std_logic                       := 'X';             -- rxblkst7
			rxsynchd0              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd0
			rxsynchd1              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd1
			rxsynchd2              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd2
			rxsynchd3              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd3
			rxsynchd4              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd4
			rxsynchd5              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd5
			rxsynchd6              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd6
			rxsynchd7              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd7
			rxfreqlocked0          : in  std_logic                       := 'X';             -- rxfreqlocked0
			rxfreqlocked1          : in  std_logic                       := 'X';             -- rxfreqlocked1
			rxfreqlocked2          : in  std_logic                       := 'X';             -- rxfreqlocked2
			rxfreqlocked3          : in  std_logic                       := 'X';             -- rxfreqlocked3
			rxfreqlocked4          : in  std_logic                       := 'X';             -- rxfreqlocked4
			rxfreqlocked5          : in  std_logic                       := 'X';             -- rxfreqlocked5
			rxfreqlocked6          : in  std_logic                       := 'X';             -- rxfreqlocked6
			rxfreqlocked7          : in  std_logic                       := 'X';             -- rxfreqlocked7
			currentcoeff0          : out std_logic_vector(17 downto 0);                      -- currentcoeff0
			currentcoeff1          : out std_logic_vector(17 downto 0);                      -- currentcoeff1
			currentcoeff2          : out std_logic_vector(17 downto 0);                      -- currentcoeff2
			currentcoeff3          : out std_logic_vector(17 downto 0);                      -- currentcoeff3
			currentcoeff4          : out std_logic_vector(17 downto 0);                      -- currentcoeff4
			currentcoeff5          : out std_logic_vector(17 downto 0);                      -- currentcoeff5
			currentcoeff6          : out std_logic_vector(17 downto 0);                      -- currentcoeff6
			currentcoeff7          : out std_logic_vector(17 downto 0);                      -- currentcoeff7
			currentrxpreset0       : out std_logic_vector(2 downto 0);                       -- currentrxpreset0
			currentrxpreset1       : out std_logic_vector(2 downto 0);                       -- currentrxpreset1
			currentrxpreset2       : out std_logic_vector(2 downto 0);                       -- currentrxpreset2
			currentrxpreset3       : out std_logic_vector(2 downto 0);                       -- currentrxpreset3
			currentrxpreset4       : out std_logic_vector(2 downto 0);                       -- currentrxpreset4
			currentrxpreset5       : out std_logic_vector(2 downto 0);                       -- currentrxpreset5
			currentrxpreset6       : out std_logic_vector(2 downto 0);                       -- currentrxpreset6
			currentrxpreset7       : out std_logic_vector(2 downto 0);                       -- currentrxpreset7
			txsynchd0              : out std_logic_vector(1 downto 0);                       -- txsynchd0
			txsynchd1              : out std_logic_vector(1 downto 0);                       -- txsynchd1
			txsynchd2              : out std_logic_vector(1 downto 0);                       -- txsynchd2
			txsynchd3              : out std_logic_vector(1 downto 0);                       -- txsynchd3
			txsynchd4              : out std_logic_vector(1 downto 0);                       -- txsynchd4
			txsynchd5              : out std_logic_vector(1 downto 0);                       -- txsynchd5
			txsynchd6              : out std_logic_vector(1 downto 0);                       -- txsynchd6
			txsynchd7              : out std_logic_vector(1 downto 0);                       -- txsynchd7
			txblkst0               : out std_logic;                                          -- txblkst0
			txblkst1               : out std_logic;                                          -- txblkst1
			txblkst2               : out std_logic;                                          -- txblkst2
			txblkst3               : out std_logic;                                          -- txblkst3
			txblkst4               : out std_logic;                                          -- txblkst4
			txblkst5               : out std_logic;                                          -- txblkst5
			txblkst6               : out std_logic;                                          -- txblkst6
			txblkst7               : out std_logic;                                          -- txblkst7
			aer_msi_num            : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- aer_msi_num
			pex_msi_num            : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- pex_msi_num
			serr_out               : out std_logic;                                          -- serr_out
			hip_reconfig_clk       : in  std_logic                       := 'X';             -- hip_reconfig_clk
			hip_reconfig_rst_n     : in  std_logic                       := 'X';             -- hip_reconfig_rst_n
			hip_reconfig_address   : in  std_logic_vector(9 downto 0)    := (others => 'X'); -- hip_reconfig_address
			hip_reconfig_read      : in  std_logic                       := 'X';             -- hip_reconfig_read
			hip_reconfig_write     : in  std_logic                       := 'X';             -- hip_reconfig_write
			hip_reconfig_writedata : in  std_logic_vector(15 downto 0)   := (others => 'X'); -- hip_reconfig_writedata
			hip_reconfig_byte_en   : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- hip_reconfig_byte_en
			ser_shift_load         : in  std_logic                       := 'X';             -- ser_shift_load
			interface_sel          : in  std_logic                       := 'X';             -- interface_sel
			cfgbp_link2csr         : in  std_logic_vector(12 downto 0)   := (others => 'X'); -- cfgbp_link2csr
			cfgbp_comclk_reg       : in  std_logic                       := 'X';             -- cfgbp_comclk_reg
			cfgbp_extsy_reg        : in  std_logic                       := 'X';             -- cfgbp_extsy_reg
			cfgbp_max_pload        : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- cfgbp_max_pload
			cfgbp_tx_ecrcgen       : in  std_logic                       := 'X';             -- cfgbp_tx_ecrcgen
			cfgbp_rx_ecrchk        : in  std_logic                       := 'X';             -- cfgbp_rx_ecrchk
			cfgbp_secbus           : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- cfgbp_secbus
			cfgbp_linkcsr_bit0     : in  std_logic                       := 'X';             -- cfgbp_linkcsr_bit0
			cfgbp_tx_req_pm        : in  std_logic                       := 'X';             -- cfgbp_tx_req_pm
			cfgbp_tx_typ_pm        : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- cfgbp_tx_typ_pm
			cfgbp_req_phypm        : in  std_logic_vector(3 downto 0)    := (others => 'X'); -- cfgbp_req_phypm
			cfgbp_req_phycfg       : in  std_logic_vector(3 downto 0)    := (others => 'X'); -- cfgbp_req_phycfg
			cfgbp_vc0_tcmap_pld    : in  std_logic_vector(6 downto 0)    := (others => 'X'); -- cfgbp_vc0_tcmap_pld
			cfgbp_inh_dllp         : in  std_logic                       := 'X';             -- cfgbp_inh_dllp
			cfgbp_inh_tx_tlp       : in  std_logic                       := 'X';             -- cfgbp_inh_tx_tlp
			cfgbp_req_wake         : in  std_logic                       := 'X';             -- cfgbp_req_wake
			cfgbp_link3_ctl        : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- cfgbp_link3_ctl
			cseb_rddata            : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- cseb_rddata
			cseb_rdresponse        : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- cseb_rdresponse
			cseb_waitrequest       : in  std_logic                       := 'X';             -- cseb_waitrequest
			cseb_wrresponse        : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- cseb_wrresponse
			cseb_wrresp_valid      : in  std_logic                       := 'X';             -- cseb_wrresp_valid
			cseb_rddata_parity     : in  std_logic_vector(3 downto 0)    := (others => 'X'); -- cseb_rddata_parity
			reservedin             : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- reservedin
			tlbfm_in               : out std_logic_vector(1000 downto 0);                    -- tlbfm_in
			tlbfm_out              : in  std_logic_vector(1000 downto 0) := (others => 'X'); -- tlbfm_out
			rxfc_cplbuf_ovf        : out std_logic                                           -- rxfc_cplbuf_ovf
		);
	end component altpcie_sv_hip_ast_hwtcl;

begin

	pcie_sv_hard_ip_inst : component altpcie_sv_hip_ast_hwtcl
		generic map (
			lane_mask_hwtcl                          => "x8",
			gen123_lane_rate_mode_hwtcl              => GEN_RATE,
			port_type_hwtcl                          => "Native endpoint",
			pcie_spec_version_hwtcl                  => "2.1",
			ast_width_hwtcl                          => "Avalon-ST 128-bit",
			pll_refclk_freq_hwtcl                    => "100 MHz",
			set_pld_clk_x1_625MHz_hwtcl              => 0,
			use_ast_parity                           => 0,
			multiple_packets_per_cycle_hwtcl         => 0,
			in_cvp_mode_hwtcl                        => 1,
			use_pci_ext_hwtcl                        => 0,
			use_pcie_ext_hwtcl                       => 0,
			use_config_bypass_hwtcl                  => 0,
			hip_reconfig_hwtcl                       => 0,
			enable_tl_only_sim_hwtcl                 => 0,
			bar0_size_mask_hwtcl                     => 13,
			bar0_io_space_hwtcl                      => "Disabled",
			bar0_64bit_mem_space_hwtcl               => "Enabled",
			bar0_prefetchable_hwtcl                  => "Enabled",
			bar1_size_mask_hwtcl                     => 0,
			bar1_io_space_hwtcl                      => "Disabled",
			bar1_prefetchable_hwtcl                  => "Disabled",
			bar2_size_mask_hwtcl                     => 13,
			bar2_io_space_hwtcl                      => "Disabled",
			bar2_64bit_mem_space_hwtcl               => "Enabled",
			bar2_prefetchable_hwtcl                  => "Enabled",
			bar3_size_mask_hwtcl                     => 0,
			bar3_io_space_hwtcl                      => "Disabled",
			bar3_prefetchable_hwtcl                  => "Disabled",
			bar4_size_mask_hwtcl                     => 22,
			bar4_io_space_hwtcl                      => "Disabled",
			bar4_64bit_mem_space_hwtcl               => "Enabled",
			bar4_prefetchable_hwtcl                  => "Enabled",
			bar5_size_mask_hwtcl                     => 0,
			bar5_io_space_hwtcl                      => "Disabled",
			bar5_prefetchable_hwtcl                  => "Disabled",
			expansion_base_address_register_hwtcl    => 0,
			io_window_addr_width_hwtcl               => 0,
			prefetchable_mem_window_addr_width_hwtcl => 0,
			vendor_id_hwtcl                          => 7103,
			device_id_hwtcl                          => DEVICE_ID,
			revision_id_hwtcl                        => 0,
			class_code_hwtcl                         => 737280,
			subsystem_vendor_id_hwtcl                => 7103,
			subsystem_device_id_hwtcl                => 7,
			max_payload_size_hwtcl                   => 128,
			extend_tag_field_hwtcl                   => "32",
			completion_timeout_hwtcl                 => "B",
			enable_completion_timeout_disable_hwtcl  => 1,
			use_aer_hwtcl                            => 1,
			ecrc_check_capable_hwtcl                 => 1,
			ecrc_gen_capable_hwtcl                   => 1,
			use_crc_forwarding_hwtcl                 => 0,
			port_link_number_hwtcl                   => 1,
			dll_active_report_support_hwtcl          => 0,
			surprise_down_error_support_hwtcl        => 0,
			slotclkcfg_hwtcl                         => 1,
			msi_multi_message_capable_hwtcl          => "4",
			msi_64bit_addressing_capable_hwtcl       => "true",
			msi_masking_capable_hwtcl                => "false",
			msi_support_hwtcl                        => "true",
			enable_function_msix_support_hwtcl       => 0,
			msix_table_size_hwtcl                    => 0,
			msix_table_offset_hwtcl                  => "0",
			msix_table_bir_hwtcl                     => 0,
			msix_pba_offset_hwtcl                    => "0",
			msix_pba_bir_hwtcl                       => 0,
			enable_slot_register_hwtcl               => 0,
			slot_power_scale_hwtcl                   => 0,
			slot_power_limit_hwtcl                   => 0,
			slot_number_hwtcl                        => 0,
			endpoint_l0_latency_hwtcl                => 0,
			endpoint_l1_latency_hwtcl                => 7,
			vsec_id_hwtcl                            => 40960,
			vsec_rev_hwtcl                           => 0,
			millisecond_cycle_count_hwtcl            => MS_CYCLE_COUNT,
			port_width_be_hwtcl                      => 16,
			port_width_data_hwtcl                    => 128,
			gen3_dcbal_en_hwtcl                      => 1,
			enable_pipe32_sim_hwtcl                  => 0,
			fixed_preset_on                          => 0,
			bypass_cdc_hwtcl                         => "false",
			enable_rx_buffer_checking_hwtcl          => "false",
			disable_link_x2_support_hwtcl            => "false",
			wrong_device_id_hwtcl                    => "disable",
			data_pack_rx_hwtcl                       => "disable",
			ltssm_1ms_timeout_hwtcl                  => "disable",
			ltssm_freqlocked_check_hwtcl             => "disable",
			deskew_comma_hwtcl                       => "skp_eieos_deskw",
			device_number_hwtcl                      => 0,
			pipex1_debug_sel_hwtcl                   => "disable",
			pclk_out_sel_hwtcl                       => "pclk",
			no_soft_reset_hwtcl                      => "false",
			maximum_current_hwtcl                    => 0,
			d1_support_hwtcl                         => "false",
			d2_support_hwtcl                         => "false",
			d0_pme_hwtcl                             => "false",
			d1_pme_hwtcl                             => "false",
			d2_pme_hwtcl                             => "false",
			d3_hot_pme_hwtcl                         => "false",
			d3_cold_pme_hwtcl                        => "false",
			low_priority_vc_hwtcl                    => "single_vc",
			disable_snoop_packet_hwtcl               => "false",
			enable_l1_aspm_hwtcl                     => "false",
			rx_ei_l0s_hwtcl                          => 0,
			enable_l0s_aspm_hwtcl                    => "false",
			aspm_config_management_hwtcl             => "true",
			l1_exit_latency_sameclock_hwtcl          => 0,
			l1_exit_latency_diffclock_hwtcl          => 0,
			hot_plug_support_hwtcl                   => 0,
			extended_tag_reset_hwtcl                 => "false",
			no_command_completed_hwtcl               => "true",
			interrupt_pin_hwtcl                      => "inta",
			bridge_port_vga_enable_hwtcl             => "false",
			bridge_port_ssid_support_hwtcl           => "false",
			ssvid_hwtcl                              => 0,
			ssid_hwtcl                               => 0,
			eie_before_nfts_count_hwtcl              => 4,
			gen2_diffclock_nfts_count_hwtcl          => 255,
			gen2_sameclock_nfts_count_hwtcl          => 255,
			l0_exit_latency_sameclock_hwtcl          => 6,
			l0_exit_latency_diffclock_hwtcl          => 6,
			atomic_op_routing_hwtcl                  => "false",
			atomic_op_completer_32bit_hwtcl          => "false",
			atomic_op_completer_64bit_hwtcl          => "false",
			cas_completer_128bit_hwtcl               => "false",
			ltr_mechanism_hwtcl                      => "false",
			tph_completer_hwtcl                      => "false",
			extended_format_field_hwtcl              => "false",
			atomic_malformed_hwtcl                   => "true",
			flr_capability_hwtcl                     => "false",
			enable_adapter_half_rate_mode_hwtcl      => "false",
			vc0_clk_enable_hwtcl                     => "true",
			register_pipe_signals_hwtcl              => "false",
			skp_os_gen3_count_hwtcl                  => 0,
			tx_cdc_almost_empty_hwtcl                => 5,
			rx_l0s_count_idl_hwtcl                   => 0,
			cdc_dummy_insert_limit_hwtcl             => 11,
			ei_delay_powerdown_count_hwtcl           => 10,
			skp_os_schedule_count_hwtcl              => 0,
			fc_init_timer_hwtcl                      => 1024,
			l01_entry_latency_hwtcl                  => 31,
			flow_control_update_count_hwtcl          => 30,
			flow_control_timeout_count_hwtcl         => 200,
			retry_buffer_last_active_address_hwtcl   => 2047,
			reserved_debug_hwtcl                     => 0,
			bypass_clk_switch_hwtcl                  => "false",
			l2_async_logic_hwtcl                     => "disable",
			indicator_hwtcl                          => 0,
			diffclock_nfts_count_hwtcl               => 128,
			sameclock_nfts_count_hwtcl               => 128,
			rx_cdc_almost_full_hwtcl                 => 12,
			tx_cdc_almost_full_hwtcl                 => 11,
			credit_buffer_allocation_aux_hwtcl       => "absolute",
			vc0_rx_flow_ctrl_posted_header_hwtcl     => 50,
			vc0_rx_flow_ctrl_posted_data_hwtcl       => 358,
			vc0_rx_flow_ctrl_nonposted_header_hwtcl  => 56,
			vc0_rx_flow_ctrl_nonposted_data_hwtcl    => 0,
			vc0_rx_flow_ctrl_compl_header_hwtcl      => 0,
			vc0_rx_flow_ctrl_compl_data_hwtcl        => 0,
			cpl_spc_header_hwtcl                     => 112,
			cpl_spc_data_hwtcl                       => 448,
			gen3_rxfreqlock_counter_hwtcl            => 0,
			gen3_skip_ph2_ph3_hwtcl                  => 0,
			g3_bypass_equlz_hwtcl                    => 0,
			cvp_data_compressed_hwtcl                => "false",
			cvp_data_encrypted_hwtcl                 => "false",
			cvp_mode_reset_hwtcl                     => "false",
			cvp_clk_reset_hwtcl                      => "false",
			cseb_cpl_status_during_cvp_hwtcl         => "completer_abort",
			core_clk_sel_hwtcl                       => "core_clk_250",
			cvp_rate_sel_hwtcl                       => "full_rate",
			g3_dis_rx_use_prst_hwtcl                 => "true",
			g3_dis_rx_use_prst_ep_hwtcl              => "true",
			deemphasis_enable_hwtcl                  => "false",
			reconfig_to_xcvr_width                   => 700,
			reconfig_from_xcvr_width                 => 460,
			single_rx_detect_hwtcl                   => 0,
			hip_hard_reset_hwtcl                     => 1,
			hwtcl_override_g2_txvod                  => 0,
			rpre_emph_a_val_hwtcl                    => 9,
			rpre_emph_b_val_hwtcl                    => 0,
			rpre_emph_c_val_hwtcl                    => 16,
			rpre_emph_d_val_hwtcl                    => 11,
			rpre_emph_e_val_hwtcl                    => 5,
			rvod_sel_a_val_hwtcl                     => 42,
			rvod_sel_b_val_hwtcl                     => 38,
			rvod_sel_c_val_hwtcl                     => 38,
			rvod_sel_d_val_hwtcl                     => 38,
			rvod_sel_e_val_hwtcl                     => 15,
			hwtcl_override_g3rxcoef                  => 0,
			gen3_coeff_1_hwtcl                       => 7,
			gen3_coeff_1_sel_hwtcl                   => "preset_1",
			gen3_coeff_1_preset_hint_hwtcl           => 0,
			gen3_coeff_1_nxtber_more_ptr_hwtcl       => 1,
			gen3_coeff_1_nxtber_more_hwtcl           => "g3_coeff_1_nxtber_more",
			gen3_coeff_1_nxtber_less_ptr_hwtcl       => 1,
			gen3_coeff_1_nxtber_less_hwtcl           => "g3_coeff_1_nxtber_less",
			gen3_coeff_1_reqber_hwtcl                => 0,
			gen3_coeff_1_ber_meas_hwtcl              => 2,
			gen3_coeff_2_hwtcl                       => 0,
			gen3_coeff_2_sel_hwtcl                   => "preset_2",
			gen3_coeff_2_preset_hint_hwtcl           => 0,
			gen3_coeff_2_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_2_nxtber_more_hwtcl           => "g3_coeff_2_nxtber_more",
			gen3_coeff_2_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_2_nxtber_less_hwtcl           => "g3_coeff_2_nxtber_less",
			gen3_coeff_2_reqber_hwtcl                => 0,
			gen3_coeff_2_ber_meas_hwtcl              => 0,
			gen3_coeff_3_hwtcl                       => 0,
			gen3_coeff_3_sel_hwtcl                   => "preset_3",
			gen3_coeff_3_preset_hint_hwtcl           => 0,
			gen3_coeff_3_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_3_nxtber_more_hwtcl           => "g3_coeff_3_nxtber_more",
			gen3_coeff_3_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_3_nxtber_less_hwtcl           => "g3_coeff_3_nxtber_less",
			gen3_coeff_3_reqber_hwtcl                => 0,
			gen3_coeff_3_ber_meas_hwtcl              => 0,
			gen3_coeff_4_hwtcl                       => 0,
			gen3_coeff_4_sel_hwtcl                   => "preset_4",
			gen3_coeff_4_preset_hint_hwtcl           => 0,
			gen3_coeff_4_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_4_nxtber_more_hwtcl           => "g3_coeff_4_nxtber_more",
			gen3_coeff_4_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_4_nxtber_less_hwtcl           => "g3_coeff_4_nxtber_less",
			gen3_coeff_4_reqber_hwtcl                => 0,
			gen3_coeff_4_ber_meas_hwtcl              => 0,
			gen3_coeff_5_hwtcl                       => 0,
			gen3_coeff_5_sel_hwtcl                   => "preset_5",
			gen3_coeff_5_preset_hint_hwtcl           => 0,
			gen3_coeff_5_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_5_nxtber_more_hwtcl           => "g3_coeff_5_nxtber_more",
			gen3_coeff_5_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_5_nxtber_less_hwtcl           => "g3_coeff_5_nxtber_less",
			gen3_coeff_5_reqber_hwtcl                => 0,
			gen3_coeff_5_ber_meas_hwtcl              => 0,
			gen3_coeff_6_hwtcl                       => 0,
			gen3_coeff_6_sel_hwtcl                   => "preset_6",
			gen3_coeff_6_preset_hint_hwtcl           => 0,
			gen3_coeff_6_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_6_nxtber_more_hwtcl           => "g3_coeff_6_nxtber_more",
			gen3_coeff_6_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_6_nxtber_less_hwtcl           => "g3_coeff_6_nxtber_less",
			gen3_coeff_6_reqber_hwtcl                => 0,
			gen3_coeff_6_ber_meas_hwtcl              => 0,
			gen3_coeff_7_hwtcl                       => 0,
			gen3_coeff_7_sel_hwtcl                   => "preset_7",
			gen3_coeff_7_preset_hint_hwtcl           => 0,
			gen3_coeff_7_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_7_nxtber_more_hwtcl           => "g3_coeff_7_nxtber_more",
			gen3_coeff_7_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_7_nxtber_less_hwtcl           => "g3_coeff_7_nxtber_less",
			gen3_coeff_7_reqber_hwtcl                => 0,
			gen3_coeff_7_ber_meas_hwtcl              => 0,
			gen3_coeff_8_hwtcl                       => 0,
			gen3_coeff_8_sel_hwtcl                   => "preset_8",
			gen3_coeff_8_preset_hint_hwtcl           => 0,
			gen3_coeff_8_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_8_nxtber_more_hwtcl           => "g3_coeff_8_nxtber_more",
			gen3_coeff_8_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_8_nxtber_less_hwtcl           => "g3_coeff_8_nxtber_less",
			gen3_coeff_8_reqber_hwtcl                => 0,
			gen3_coeff_8_ber_meas_hwtcl              => 0,
			gen3_coeff_9_hwtcl                       => 0,
			gen3_coeff_9_sel_hwtcl                   => "preset_9",
			gen3_coeff_9_preset_hint_hwtcl           => 0,
			gen3_coeff_9_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_9_nxtber_more_hwtcl           => "g3_coeff_9_nxtber_more",
			gen3_coeff_9_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_9_nxtber_less_hwtcl           => "g3_coeff_9_nxtber_less",
			gen3_coeff_9_reqber_hwtcl                => 0,
			gen3_coeff_9_ber_meas_hwtcl              => 0,
			gen3_coeff_10_hwtcl                      => 0,
			gen3_coeff_10_sel_hwtcl                  => "preset_10",
			gen3_coeff_10_preset_hint_hwtcl          => 0,
			gen3_coeff_10_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_10_nxtber_more_hwtcl          => "g3_coeff_10_nxtber_more",
			gen3_coeff_10_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_10_nxtber_less_hwtcl          => "g3_coeff_10_nxtber_less",
			gen3_coeff_10_reqber_hwtcl               => 0,
			gen3_coeff_10_ber_meas_hwtcl             => 0,
			gen3_coeff_11_hwtcl                      => 0,
			gen3_coeff_11_sel_hwtcl                  => "preset_11",
			gen3_coeff_11_preset_hint_hwtcl          => 0,
			gen3_coeff_11_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_11_nxtber_more_hwtcl          => "g3_coeff_11_nxtber_more",
			gen3_coeff_11_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_11_nxtber_less_hwtcl          => "g3_coeff_11_nxtber_less",
			gen3_coeff_11_reqber_hwtcl               => 0,
			gen3_coeff_11_ber_meas_hwtcl             => 0,
			gen3_coeff_12_hwtcl                      => 0,
			gen3_coeff_12_sel_hwtcl                  => "preset_12",
			gen3_coeff_12_preset_hint_hwtcl          => 0,
			gen3_coeff_12_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_12_nxtber_more_hwtcl          => "g3_coeff_12_nxtber_more",
			gen3_coeff_12_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_12_nxtber_less_hwtcl          => "g3_coeff_12_nxtber_less",
			gen3_coeff_12_reqber_hwtcl               => 0,
			gen3_coeff_12_ber_meas_hwtcl             => 0,
			gen3_coeff_13_hwtcl                      => 0,
			gen3_coeff_13_sel_hwtcl                  => "preset_13",
			gen3_coeff_13_preset_hint_hwtcl          => 0,
			gen3_coeff_13_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_13_nxtber_more_hwtcl          => "g3_coeff_13_nxtber_more",
			gen3_coeff_13_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_13_nxtber_less_hwtcl          => "g3_coeff_13_nxtber_less",
			gen3_coeff_13_reqber_hwtcl               => 0,
			gen3_coeff_13_ber_meas_hwtcl             => 0,
			gen3_coeff_14_hwtcl                      => 0,
			gen3_coeff_14_sel_hwtcl                  => "preset_14",
			gen3_coeff_14_preset_hint_hwtcl          => 0,
			gen3_coeff_14_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_14_nxtber_more_hwtcl          => "g3_coeff_14_nxtber_more",
			gen3_coeff_14_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_14_nxtber_less_hwtcl          => "g3_coeff_14_nxtber_less",
			gen3_coeff_14_reqber_hwtcl               => 0,
			gen3_coeff_14_ber_meas_hwtcl             => 0,
			gen3_coeff_15_hwtcl                      => 0,
			gen3_coeff_15_sel_hwtcl                  => "preset_15",
			gen3_coeff_15_preset_hint_hwtcl          => 0,
			gen3_coeff_15_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_15_nxtber_more_hwtcl          => "g3_coeff_15_nxtber_more",
			gen3_coeff_15_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_15_nxtber_less_hwtcl          => "g3_coeff_15_nxtber_less",
			gen3_coeff_15_reqber_hwtcl               => 0,
			gen3_coeff_15_ber_meas_hwtcl             => 0,
			gen3_coeff_16_hwtcl                      => 0,
			gen3_coeff_16_sel_hwtcl                  => "preset_16",
			gen3_coeff_16_preset_hint_hwtcl          => 0,
			gen3_coeff_16_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_16_nxtber_more_hwtcl          => "g3_coeff_16_nxtber_more",
			gen3_coeff_16_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_16_nxtber_less_hwtcl          => "g3_coeff_16_nxtber_less",
			gen3_coeff_16_reqber_hwtcl               => 0,
			gen3_coeff_16_ber_meas_hwtcl             => 0,
			gen3_coeff_17_hwtcl                      => 0,
			gen3_coeff_17_sel_hwtcl                  => "preset_17",
			gen3_coeff_17_preset_hint_hwtcl          => 0,
			gen3_coeff_17_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_17_nxtber_more_hwtcl          => "g3_coeff_17_nxtber_more",
			gen3_coeff_17_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_17_nxtber_less_hwtcl          => "g3_coeff_17_nxtber_less",
			gen3_coeff_17_reqber_hwtcl               => 0,
			gen3_coeff_17_ber_meas_hwtcl             => 0,
			gen3_coeff_18_hwtcl                      => 0,
			gen3_coeff_18_sel_hwtcl                  => "preset_18",
			gen3_coeff_18_preset_hint_hwtcl          => 0,
			gen3_coeff_18_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_18_nxtber_more_hwtcl          => "g3_coeff_18_nxtber_more",
			gen3_coeff_18_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_18_nxtber_less_hwtcl          => "g3_coeff_18_nxtber_less",
			gen3_coeff_18_reqber_hwtcl               => 0,
			gen3_coeff_18_ber_meas_hwtcl             => 0,
			gen3_coeff_19_hwtcl                      => 0,
			gen3_coeff_19_sel_hwtcl                  => "preset_19",
			gen3_coeff_19_preset_hint_hwtcl          => 0,
			gen3_coeff_19_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_19_nxtber_more_hwtcl          => "g3_coeff_19_nxtber_more",
			gen3_coeff_19_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_19_nxtber_less_hwtcl          => "g3_coeff_19_nxtber_less",
			gen3_coeff_19_reqber_hwtcl               => 0,
			gen3_coeff_19_ber_meas_hwtcl             => 0,
			gen3_coeff_20_hwtcl                      => 0,
			gen3_coeff_20_sel_hwtcl                  => "preset_20",
			gen3_coeff_20_preset_hint_hwtcl          => 0,
			gen3_coeff_20_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_20_nxtber_more_hwtcl          => "g3_coeff_20_nxtber_more",
			gen3_coeff_20_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_20_nxtber_less_hwtcl          => "g3_coeff_20_nxtber_less",
			gen3_coeff_20_reqber_hwtcl               => 0,
			gen3_coeff_20_ber_meas_hwtcl             => 0,
			gen3_coeff_21_hwtcl                      => 0,
			gen3_coeff_21_sel_hwtcl                  => "preset_21",
			gen3_coeff_21_preset_hint_hwtcl          => 0,
			gen3_coeff_21_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_21_nxtber_more_hwtcl          => "g3_coeff_21_nxtber_more",
			gen3_coeff_21_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_21_nxtber_less_hwtcl          => "g3_coeff_21_nxtber_less",
			gen3_coeff_21_reqber_hwtcl               => 0,
			gen3_coeff_21_ber_meas_hwtcl             => 0,
			gen3_coeff_22_hwtcl                      => 0,
			gen3_coeff_22_sel_hwtcl                  => "preset_22",
			gen3_coeff_22_preset_hint_hwtcl          => 0,
			gen3_coeff_22_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_22_nxtber_more_hwtcl          => "g3_coeff_22_nxtber_more",
			gen3_coeff_22_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_22_nxtber_less_hwtcl          => "g3_coeff_22_nxtber_less",
			gen3_coeff_22_reqber_hwtcl               => 0,
			gen3_coeff_22_ber_meas_hwtcl             => 0,
			gen3_coeff_23_hwtcl                      => 0,
			gen3_coeff_23_sel_hwtcl                  => "preset_23",
			gen3_coeff_23_preset_hint_hwtcl          => 0,
			gen3_coeff_23_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_23_nxtber_more_hwtcl          => "g3_coeff_23_nxtber_more",
			gen3_coeff_23_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_23_nxtber_less_hwtcl          => "g3_coeff_23_nxtber_less",
			gen3_coeff_23_reqber_hwtcl               => 0,
			gen3_coeff_23_ber_meas_hwtcl             => 0,
			gen3_coeff_24_hwtcl                      => 0,
			gen3_coeff_24_sel_hwtcl                  => "preset_24",
			gen3_coeff_24_preset_hint_hwtcl          => 0,
			gen3_coeff_24_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_24_nxtber_more_hwtcl          => "g3_coeff_24_nxtber_more",
			gen3_coeff_24_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_24_nxtber_less_hwtcl          => "g3_coeff_24_nxtber_less",
			gen3_coeff_24_reqber_hwtcl               => 0,
			gen3_coeff_24_ber_meas_hwtcl             => 0,
			hwtcl_override_g3txcoef                  => 0,
			gen3_preset_coeff_1_hwtcl                => 0,
			gen3_preset_coeff_2_hwtcl                => 0,
			gen3_preset_coeff_3_hwtcl                => 0,
			gen3_preset_coeff_4_hwtcl                => 0,
			gen3_preset_coeff_5_hwtcl                => 0,
			gen3_preset_coeff_6_hwtcl                => 0,
			gen3_preset_coeff_7_hwtcl                => 0,
			gen3_preset_coeff_8_hwtcl                => 0,
			gen3_preset_coeff_9_hwtcl                => 0,
			gen3_preset_coeff_10_hwtcl               => 0,
			gen3_preset_coeff_11_hwtcl               => 0,
			gen3_low_freq_hwtcl                      => 0,
			full_swing_hwtcl                         => 53,
			gen3_full_swing_hwtcl                    => 35,
			use_atx_pll_hwtcl                        => 0,
			low_latency_mode_hwtcl                   => 0
		)
		port map (
			npor                   => npor,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --               npor.npor
			pin_perst              => pin_perst,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .pin_perst
			lmi_addr               => lmi_addr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                lmi.lmi_addr
			lmi_din                => lmi_din,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .lmi_din
			lmi_rden               => lmi_rden,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .lmi_rden
			lmi_wren               => lmi_wren,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .lmi_wren
			lmi_ack                => lmi_ack,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .lmi_ack
			lmi_dout               => lmi_dout,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .lmi_dout
			hpg_ctrler             => hpg_ctrler,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --          config_tl.hpg_ctrler
			tl_cfg_add             => tl_cfg_add,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .tl_cfg_add
			tl_cfg_ctl             => tl_cfg_ctl,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .tl_cfg_ctl
			tl_cfg_sts             => tl_cfg_sts,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .tl_cfg_sts
			cpl_err                => cpl_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .cpl_err
			cpl_pending            => cpl_pending,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .cpl_pending
			pm_auxpwr              => pm_auxpwr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --         power_mngt.pm_auxpwr
			pm_data                => pm_data,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .pm_data
			pme_to_cr              => pme_to_cr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .pme_to_cr
			pm_event               => pm_event,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .pm_event
			pme_to_sr              => pme_to_sr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .pme_to_sr
			rx_st_sop              => rx_st_sop,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --              rx_st.startofpacket
			rx_st_eop              => rx_st_eop,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .endofpacket
			rx_st_err              => rx_st_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .error
			rx_st_valid            => rx_st_valid,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .valid
			rx_st_empty            => rx_st_empty,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .empty
			rx_st_ready            => rx_st_ready,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .ready
			rx_st_data             => rx_st_data,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .data
			rx_st_bar              => rx_st_bar,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --          rx_bar_be.rx_st_bar
			rx_st_mask             => rx_st_mask,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .rx_st_mask
			tx_st_sop              => tx_st_sop,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --              tx_st.startofpacket
			tx_st_eop              => tx_st_eop,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .endofpacket
			tx_st_err              => tx_st_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .error
			tx_st_valid            => tx_st_valid,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .valid
			tx_st_empty            => tx_st_empty,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .empty
			tx_st_ready            => tx_st_ready,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .ready
			tx_st_data             => tx_st_data,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .data
			tx_cred_datafccp       => tx_cred_datafccp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --            tx_cred.tx_cred_datafccp
			tx_cred_datafcnp       => tx_cred_datafcnp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .tx_cred_datafcnp
			tx_cred_datafcp        => tx_cred_datafcp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .tx_cred_datafcp
			tx_cred_fchipcons      => tx_cred_fchipcons,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .tx_cred_fchipcons
			tx_cred_fcinfinite     => tx_cred_fcinfinite,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .tx_cred_fcinfinite
			tx_cred_hdrfccp        => tx_cred_hdrfccp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .tx_cred_hdrfccp
			tx_cred_hdrfcnp        => tx_cred_hdrfcnp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .tx_cred_hdrfcnp
			tx_cred_hdrfcp         => tx_cred_hdrfcp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_cred_hdrfcp
			pld_clk                => pld_clk,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --            pld_clk.clk
			coreclkout_hip         => coreclkout_hip,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --     coreclkout_hip.clk
			refclk                 => refclk,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --             refclk.clk
			reset_status           => reset_status,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --            hip_rst.reset_status
			serdes_pll_locked      => serdes_pll_locked,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .serdes_pll_locked
			pld_clk_inuse          => pld_clk_inuse,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --                   .pld_clk_inuse
			pld_core_ready         => pld_core_ready,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .pld_core_ready
			testin_zero            => testin_zero,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .testin_zero
			reconfig_to_xcvr       => reconfig_to_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr     => reconfig_from_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          -- reconfig_from_xcvr.reconfig_from_xcvr
			rx_in0                 => rx_in0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --         hip_serial.rx_in0
			rx_in1                 => rx_in1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .rx_in1
			rx_in2                 => rx_in2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .rx_in2
			rx_in3                 => rx_in3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .rx_in3
			rx_in4                 => rx_in4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .rx_in4
			rx_in5                 => rx_in5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .rx_in5
			rx_in6                 => rx_in6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .rx_in6
			rx_in7                 => rx_in7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .rx_in7
			tx_out0                => tx_out0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .tx_out0
			tx_out1                => tx_out1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .tx_out1
			tx_out2                => tx_out2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .tx_out2
			tx_out3                => tx_out3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .tx_out3
			tx_out4                => tx_out4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .tx_out4
			tx_out5                => tx_out5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .tx_out5
			tx_out6                => tx_out6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .tx_out6
			tx_out7                => tx_out7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .tx_out7
			sim_pipe_pclk_in       => sim_pipe_pclk_in,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --           hip_pipe.sim_pipe_pclk_in
			sim_pipe_rate          => sim_pipe_rate,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --                   .sim_pipe_rate
			sim_ltssmstate         => sim_ltssmstate,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .sim_ltssmstate
			eidleinfersel0         => eidleinfersel0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .eidleinfersel0
			eidleinfersel1         => eidleinfersel1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .eidleinfersel1
			eidleinfersel2         => eidleinfersel2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .eidleinfersel2
			eidleinfersel3         => eidleinfersel3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .eidleinfersel3
			eidleinfersel4         => eidleinfersel4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .eidleinfersel4
			eidleinfersel5         => eidleinfersel5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .eidleinfersel5
			eidleinfersel6         => eidleinfersel6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .eidleinfersel6
			eidleinfersel7         => eidleinfersel7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .eidleinfersel7
			powerdown0             => powerdown0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .powerdown0
			powerdown1             => powerdown1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .powerdown1
			powerdown2             => powerdown2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .powerdown2
			powerdown3             => powerdown3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .powerdown3
			powerdown4             => powerdown4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .powerdown4
			powerdown5             => powerdown5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .powerdown5
			powerdown6             => powerdown6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .powerdown6
			powerdown7             => powerdown7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .powerdown7
			rxpolarity0            => rxpolarity0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxpolarity0
			rxpolarity1            => rxpolarity1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxpolarity1
			rxpolarity2            => rxpolarity2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxpolarity2
			rxpolarity3            => rxpolarity3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxpolarity3
			rxpolarity4            => rxpolarity4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxpolarity4
			rxpolarity5            => rxpolarity5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxpolarity5
			rxpolarity6            => rxpolarity6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxpolarity6
			rxpolarity7            => rxpolarity7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxpolarity7
			txcompl0               => txcompl0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txcompl0
			txcompl1               => txcompl1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txcompl1
			txcompl2               => txcompl2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txcompl2
			txcompl3               => txcompl3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txcompl3
			txcompl4               => txcompl4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txcompl4
			txcompl5               => txcompl5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txcompl5
			txcompl6               => txcompl6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txcompl6
			txcompl7               => txcompl7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txcompl7
			txdata0                => txdata0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .txdata0
			txdata1                => txdata1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .txdata1
			txdata2                => txdata2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .txdata2
			txdata3                => txdata3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .txdata3
			txdata4                => txdata4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .txdata4
			txdata5                => txdata5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .txdata5
			txdata6                => txdata6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .txdata6
			txdata7                => txdata7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .txdata7
			txdatak0               => txdatak0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txdatak0
			txdatak1               => txdatak1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txdatak1
			txdatak2               => txdatak2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txdatak2
			txdatak3               => txdatak3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txdatak3
			txdatak4               => txdatak4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txdatak4
			txdatak5               => txdatak5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txdatak5
			txdatak6               => txdatak6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txdatak6
			txdatak7               => txdatak7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txdatak7
			txdetectrx0            => txdetectrx0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txdetectrx0
			txdetectrx1            => txdetectrx1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txdetectrx1
			txdetectrx2            => txdetectrx2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txdetectrx2
			txdetectrx3            => txdetectrx3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txdetectrx3
			txdetectrx4            => txdetectrx4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txdetectrx4
			txdetectrx5            => txdetectrx5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txdetectrx5
			txdetectrx6            => txdetectrx6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txdetectrx6
			txdetectrx7            => txdetectrx7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txdetectrx7
			txelecidle0            => txelecidle0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txelecidle0
			txelecidle1            => txelecidle1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txelecidle1
			txelecidle2            => txelecidle2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txelecidle2
			txelecidle3            => txelecidle3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txelecidle3
			txelecidle4            => txelecidle4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txelecidle4
			txelecidle5            => txelecidle5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txelecidle5
			txelecidle6            => txelecidle6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txelecidle6
			txelecidle7            => txelecidle7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .txelecidle7
			txdeemph0              => txdeemph0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txdeemph0
			txdeemph1              => txdeemph1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txdeemph1
			txdeemph2              => txdeemph2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txdeemph2
			txdeemph3              => txdeemph3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txdeemph3
			txdeemph4              => txdeemph4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txdeemph4
			txdeemph5              => txdeemph5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txdeemph5
			txdeemph6              => txdeemph6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txdeemph6
			txdeemph7              => txdeemph7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txdeemph7
			txmargin0              => txmargin0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txmargin0
			txmargin1              => txmargin1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txmargin1
			txmargin2              => txmargin2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txmargin2
			txmargin3              => txmargin3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txmargin3
			txmargin4              => txmargin4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txmargin4
			txmargin5              => txmargin5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txmargin5
			txmargin6              => txmargin6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txmargin6
			txmargin7              => txmargin7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .txmargin7
			txswing0               => txswing0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txswing0
			txswing1               => txswing1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txswing1
			txswing2               => txswing2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txswing2
			txswing3               => txswing3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txswing3
			txswing4               => txswing4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txswing4
			txswing5               => txswing5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txswing5
			txswing6               => txswing6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txswing6
			txswing7               => txswing7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .txswing7
			phystatus0             => phystatus0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .phystatus0
			phystatus1             => phystatus1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .phystatus1
			phystatus2             => phystatus2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .phystatus2
			phystatus3             => phystatus3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .phystatus3
			phystatus4             => phystatus4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .phystatus4
			phystatus5             => phystatus5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .phystatus5
			phystatus6             => phystatus6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .phystatus6
			phystatus7             => phystatus7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .phystatus7
			rxdata0                => rxdata0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .rxdata0
			rxdata1                => rxdata1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .rxdata1
			rxdata2                => rxdata2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .rxdata2
			rxdata3                => rxdata3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .rxdata3
			rxdata4                => rxdata4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .rxdata4
			rxdata5                => rxdata5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .rxdata5
			rxdata6                => rxdata6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .rxdata6
			rxdata7                => rxdata7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .rxdata7
			rxdatak0               => rxdatak0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxdatak0
			rxdatak1               => rxdatak1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxdatak1
			rxdatak2               => rxdatak2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxdatak2
			rxdatak3               => rxdatak3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxdatak3
			rxdatak4               => rxdatak4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxdatak4
			rxdatak5               => rxdatak5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxdatak5
			rxdatak6               => rxdatak6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxdatak6
			rxdatak7               => rxdatak7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxdatak7
			rxelecidle0            => rxelecidle0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxelecidle0
			rxelecidle1            => rxelecidle1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxelecidle1
			rxelecidle2            => rxelecidle2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxelecidle2
			rxelecidle3            => rxelecidle3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxelecidle3
			rxelecidle4            => rxelecidle4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxelecidle4
			rxelecidle5            => rxelecidle5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxelecidle5
			rxelecidle6            => rxelecidle6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxelecidle6
			rxelecidle7            => rxelecidle7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .rxelecidle7
			rxstatus0              => rxstatus0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .rxstatus0
			rxstatus1              => rxstatus1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .rxstatus1
			rxstatus2              => rxstatus2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .rxstatus2
			rxstatus3              => rxstatus3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .rxstatus3
			rxstatus4              => rxstatus4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .rxstatus4
			rxstatus5              => rxstatus5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .rxstatus5
			rxstatus6              => rxstatus6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .rxstatus6
			rxstatus7              => rxstatus7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .rxstatus7
			rxvalid0               => rxvalid0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxvalid0
			rxvalid1               => rxvalid1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxvalid1
			rxvalid2               => rxvalid2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxvalid2
			rxvalid3               => rxvalid3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxvalid3
			rxvalid4               => rxvalid4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxvalid4
			rxvalid5               => rxvalid5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxvalid5
			rxvalid6               => rxvalid6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxvalid6
			rxvalid7               => rxvalid7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rxvalid7
			app_int_sts            => app_int_sts,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --            int_msi.app_int_sts
			app_msi_num            => app_msi_num,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .app_msi_num
			app_msi_req            => app_msi_req,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .app_msi_req
			app_msi_tc             => app_msi_tc,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .app_msi_tc
			app_int_ack            => app_int_ack,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .app_int_ack
			app_msi_ack            => app_msi_ack,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .app_msi_ack
			test_in                => test_in,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --           hip_ctrl.test_in
			simu_mode_pipe         => simu_mode_pipe,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .simu_mode_pipe
			derr_cor_ext_rcv       => derr_cor_ext_rcv,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --         hip_status.derr_cor_ext_rcv
			derr_cor_ext_rpl       => derr_cor_ext_rpl,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .derr_cor_ext_rpl
			derr_rpl               => derr_rpl,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .derr_rpl
			dlup                   => dlup,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .dlup
			dlup_exit              => dlup_exit,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .dlup_exit
			ev128ns                => ev128ns,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .ev128ns
			ev1us                  => ev1us,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --                   .ev1us
			hotrst_exit            => hotrst_exit,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .hotrst_exit
			int_status             => int_status,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .int_status
			l2_exit                => l2_exit,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .l2_exit
			lane_act               => lane_act,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .lane_act
			ltssmstate             => ltssmstate,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .ltssmstate
			rx_par_err             => rx_par_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .rx_par_err
			tx_par_err             => tx_par_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .tx_par_err
			cfg_par_err            => cfg_par_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .cfg_par_err
			ko_cpl_spc_header      => ko_cpl_spc_header,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .ko_cpl_spc_header
			ko_cpl_spc_data        => ko_cpl_spc_data,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .ko_cpl_spc_data
			currentspeed           => currentspeed,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --   hip_currentspeed.currentspeed
			rx_st_parity           => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rx_st_be               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			tx_st_parity           => "0000000000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --        (terminated)
			tx_cons_cred_sel       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			sim_pipe_pclk_out      => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxdataskip0            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip1            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip2            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip3            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip4            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip5            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip6            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip7            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst0               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst1               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst2               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst3               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst4               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst5               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst6               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst7               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxsynchd0              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd1              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd2              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd3              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd4              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd5              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd6              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd7              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxfreqlocked0          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked1          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked2          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked3          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked4          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked5          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked6          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked7          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			currentcoeff0          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff1          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff2          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff3          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff4          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff5          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff6          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff7          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset0       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset1       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset2       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset3       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset4       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset5       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset6       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset7       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd0              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd1              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd2              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd3              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd4              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd5              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd6              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd7              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst0               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst1               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst2               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst3               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst4               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst5               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst6               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst7               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			aer_msi_num            => "00000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --        (terminated)
			pex_msi_num            => "00000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --        (terminated)
			serr_out               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			hip_reconfig_clk       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			hip_reconfig_rst_n     => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			hip_reconfig_address   => "0000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			hip_reconfig_read      => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			hip_reconfig_write     => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			hip_reconfig_writedata => "0000000000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --        (terminated)
			hip_reconfig_byte_en   => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			ser_shift_load         => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			interface_sel          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_link2csr         => "0000000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --        (terminated)
			cfgbp_comclk_reg       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_extsy_reg        => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_max_pload        => "000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --        (terminated)
			cfgbp_tx_ecrcgen       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_rx_ecrchk        => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_secbus           => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --        (terminated)
			cfgbp_linkcsr_bit0     => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_tx_req_pm        => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_tx_typ_pm        => "000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --        (terminated)
			cfgbp_req_phypm        => "0000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --        (terminated)
			cfgbp_req_phycfg       => "0000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --        (terminated)
			cfgbp_vc0_tcmap_pld    => "0000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --        (terminated)
			cfgbp_inh_dllp         => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_inh_tx_tlp       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_req_wake         => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_link3_ctl        => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			cseb_rddata            => "00000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --        (terminated)
			cseb_rdresponse        => "00000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --        (terminated)
			cseb_waitrequest       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cseb_wrresponse        => "00000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --        (terminated)
			cseb_wrresp_valid      => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cseb_rddata_parity     => "0000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --        (terminated)
			reservedin             => "00000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --        (terminated)
			tlbfm_in               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			tlbfm_out              => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			rxfc_cplbuf_ovf        => open                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
		);

end architecture rtl; -- of pcie_SV_hard_ip
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2013 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_pcie_sv_hip_ast" version="13.1" >
-- Retrieval info: 	<generic name="design_environment_hwtcl" value="NATIVE" />
-- Retrieval info: 	<generic name="INTENDED_DEVICE_FAMILY" value="Stratix" />
-- Retrieval info: 	<generic name="pcie_qsys" value="1" />
-- Retrieval info: 	<generic name="lane_mask_hwtcl" value="x8" />
-- Retrieval info: 	<generic name="gen123_lane_rate_mode_hwtcl" value="Gen2 (5.0 Gbps)" />
-- Retrieval info: 	<generic name="port_type_hwtcl" value="Native endpoint" />
-- Retrieval info: 	<generic name="pcie_spec_version_hwtcl" value="2.1" />
-- Retrieval info: 	<generic name="ast_width_hwtcl" value="Avalon-ST 128-bit" />
-- Retrieval info: 	<generic name="rxbuffer_rxreq_hwtcl" value="Balanced" />
-- Retrieval info: 	<generic name="pll_refclk_freq_hwtcl" value="100 MHz" />
-- Retrieval info: 	<generic name="set_pld_clk_x1_625MHz_hwtcl" value="0" />
-- Retrieval info: 	<generic name="use_rx_st_be_hwtcl" value="0" />
-- Retrieval info: 	<generic name="use_ast_parity" value="0" />
-- Retrieval info: 	<generic name="multiple_packets_per_cycle_hwtcl" value="0" />
-- Retrieval info: 	<generic name="in_cvp_mode_hwtcl" value="1" />
-- Retrieval info: 	<generic name="use_tx_cons_cred_sel_hwtcl" value="0" />
-- Retrieval info: 	<generic name="use_pci_ext_hwtcl" value="0" />
-- Retrieval info: 	<generic name="use_pcie_ext_hwtcl" value="0" />
-- Retrieval info: 	<generic name="use_config_bypass_hwtcl" value="0" />
-- Retrieval info: 	<generic name="hip_reconfig_hwtcl" value="0" />
-- Retrieval info: 	<generic name="enable_tl_only_sim_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar0_type_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar0_size_mask_hwtcl" value="13" />
-- Retrieval info: 	<generic name="bar1_type_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar1_size_mask_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_type_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar2_size_mask_hwtcl" value="13" />
-- Retrieval info: 	<generic name="bar3_type_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_size_mask_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_type_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar4_size_mask_hwtcl" value="22" />
-- Retrieval info: 	<generic name="bar5_type_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_size_mask_hwtcl" value="0" />
-- Retrieval info: 	<generic name="expansion_base_address_register_hwtcl" value="0" />
-- Retrieval info: 	<generic name="io_window_addr_width_hwtcl" value="0" />
-- Retrieval info: 	<generic name="prefetchable_mem_window_addr_width_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vendor_id_hwtcl" value="7103" />
-- Retrieval info: 	<generic name="device_id_hwtcl" value="4" />
-- Retrieval info: 	<generic name="revision_id_hwtcl" value="0" />
-- Retrieval info: 	<generic name="class_code_hwtcl" value="737280" />
-- Retrieval info: 	<generic name="subsystem_vendor_id_hwtcl" value="7103" />
-- Retrieval info: 	<generic name="subsystem_device_id_hwtcl" value="7" />
-- Retrieval info: 	<generic name="max_payload_size_hwtcl" value="128" />
-- Retrieval info: 	<generic name="extend_tag_field_hwtcl" value="32" />
-- Retrieval info: 	<generic name="completion_timeout_hwtcl" value="B" />
-- Retrieval info: 	<generic name="enable_completion_timeout_disable_hwtcl" value="1" />
-- Retrieval info: 	<generic name="use_aer_hwtcl" value="1" />
-- Retrieval info: 	<generic name="ecrc_check_capable_hwtcl" value="1" />
-- Retrieval info: 	<generic name="ecrc_gen_capable_hwtcl" value="1" />
-- Retrieval info: 	<generic name="use_crc_forwarding_hwtcl" value="0" />
-- Retrieval info: 	<generic name="track_rxfc_cplbuf_ovf_hwtcl" value="0" />
-- Retrieval info: 	<generic name="port_link_number_hwtcl" value="1" />
-- Retrieval info: 	<generic name="dll_active_report_support_hwtcl" value="0" />
-- Retrieval info: 	<generic name="surprise_down_error_support_hwtcl" value="0" />
-- Retrieval info: 	<generic name="slotclkcfg_hwtcl" value="1" />
-- Retrieval info: 	<generic name="msi_multi_message_capable_hwtcl" value="4" />
-- Retrieval info: 	<generic name="msi_64bit_addressing_capable_hwtcl" value="true" />
-- Retrieval info: 	<generic name="msi_masking_capable_hwtcl" value="false" />
-- Retrieval info: 	<generic name="msi_support_hwtcl" value="true" />
-- Retrieval info: 	<generic name="enable_function_msix_support_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_size_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_offset_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_bir_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_offset_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_bir_hwtcl" value="0" />
-- Retrieval info: 	<generic name="enable_slot_register_hwtcl" value="0" />
-- Retrieval info: 	<generic name="slot_power_scale_hwtcl" value="0" />
-- Retrieval info: 	<generic name="slot_power_limit_hwtcl" value="0" />
-- Retrieval info: 	<generic name="slot_number_hwtcl" value="0" />
-- Retrieval info: 	<generic name="endpoint_l0_latency_hwtcl" value="0" />
-- Retrieval info: 	<generic name="endpoint_l1_latency_hwtcl" value="7" />
-- Retrieval info: 	<generic name="vsec_id_hwtcl" value="40960" />
-- Retrieval info: 	<generic name="vsec_rev_hwtcl" value="0" />
-- Retrieval info: 	<generic name="enable_pipe32_sim_hwtcl" value="0" />
-- Retrieval info: 	<generic name="enable_pipe32_phyip_ser_driver_hwtcl" value="0" />
-- Retrieval info: 	<generic name="fixed_preset_on" value="0" />
-- Retrieval info: 	<generic name="advanced_default_parameter_override" value="0" />
-- Retrieval info: 	<generic name="override_tbpartner_driver_setting_hwtcl" value="0" />
-- Retrieval info: 	<generic name="override_rxbuffer_cred_preset" value="0" />
-- Retrieval info: 	<generic name="gen3_rxfreqlock_counter_hwtcl" value="0" />
-- Retrieval info: 	<generic name="force_hrc" value="0" />
-- Retrieval info: 	<generic name="force_src" value="0" />
-- Retrieval info: 	<generic name="serial_sim_hwtcl" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_bypass_cdc" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_enable_rx_buffer_checking" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_disable_link_x2_support" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_wrong_device_id" value="disable" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_data_pack_rx" value="disable" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_ltssm_1ms_timeout" value="disable" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_ltssm_freqlocked_check" value="disable" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_deskew_comma" value="com_deskw" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_device_number" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_pipex1_debug_sel" value="disable" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_pclk_out_sel" value="pclk" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_no_soft_reset" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_maximum_current" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_d1_support" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_d2_support" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_d0_pme" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_d1_pme" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_d2_pme" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_d3_hot_pme" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_d3_cold_pme" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_low_priority_vc" value="single_vc" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_disable_snoop_packet" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_enable_l1_aspm" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_set_l0s" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_l1_exit_latency_sameclock" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_l1_exit_latency_diffclock" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_hot_plug_support" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_extended_tag_reset" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_no_command_completed" value="true" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_interrupt_pin" value="inta" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_bridge_port_vga_enable" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_bridge_port_ssid_support" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_ssvid" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_ssid" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_eie_before_nfts_count" value="4" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_gen2_diffclock_nfts_count" value="255" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_gen2_sameclock_nfts_count" value="255" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_l0_exit_latency_sameclock" value="6" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_l0_exit_latency_diffclock" value="6" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_atomic_op_routing" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_atomic_op_completer_32bit" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_atomic_op_completer_64bit" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_cas_completer_128bit" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_ltr_mechanism" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_tph_completer" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_extended_format_field" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_atomic_malformed" value="true" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_flr_capability" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_enable_adapter_half_rate_mode" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_vc0_clk_enable" value="true" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_register_pipe_signals" value="false" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_skp_os_gen3_count" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_tx_cdc_almost_empty" value="5" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_rx_l0s_count_idl" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_cdc_dummy_insert_limit" value="11" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_ei_delay_powerdown_count" value="10" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_skp_os_schedule_count" value="0" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_fc_init_timer" value="1024" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_l01_entry_latency" value="31" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_flow_control_update_count" value="30" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_flow_control_timeout_count" value="200" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_retry_buffer_last_active_address" value="2047" />
-- Retrieval info: 	<generic name="advanced_default_hwtcl_reserved_debug" value="0" />
-- Retrieval info: 	<generic name="hwtcl_override_g2_txvod" value="0" />
-- Retrieval info: 	<generic name="rpre_emph_a_val_hwtcl" value="9" />
-- Retrieval info: 	<generic name="rpre_emph_b_val_hwtcl" value="0" />
-- Retrieval info: 	<generic name="rpre_emph_c_val_hwtcl" value="16" />
-- Retrieval info: 	<generic name="rpre_emph_d_val_hwtcl" value="11" />
-- Retrieval info: 	<generic name="rpre_emph_e_val_hwtcl" value="5" />
-- Retrieval info: 	<generic name="rvod_sel_a_val_hwtcl" value="42" />
-- Retrieval info: 	<generic name="rvod_sel_b_val_hwtcl" value="38" />
-- Retrieval info: 	<generic name="rvod_sel_c_val_hwtcl" value="38" />
-- Retrieval info: 	<generic name="rvod_sel_d_val_hwtcl" value="38" />
-- Retrieval info: 	<generic name="rvod_sel_e_val_hwtcl" value="15" />
-- Retrieval info: 	<generic name="hwtcl_override_g3rxcoef" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_1_hwtcl" value="7" />
-- Retrieval info: 	<generic name="gen3_coeff_1_sel_hwtcl" value="preset_1" />
-- Retrieval info: 	<generic name="gen3_coeff_1_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_1_nxtber_more_ptr_hwtcl" value="1" />
-- Retrieval info: 	<generic name="gen3_coeff_1_nxtber_more_hwtcl" value="g3_coeff_1_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_1_nxtber_less_ptr_hwtcl" value="1" />
-- Retrieval info: 	<generic name="gen3_coeff_1_nxtber_less_hwtcl" value="g3_coeff_1_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_1_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_1_ber_meas_hwtcl" value="2" />
-- Retrieval info: 	<generic name="gen3_coeff_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_2_sel_hwtcl" value="preset_2" />
-- Retrieval info: 	<generic name="gen3_coeff_2_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_2_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_2_nxtber_more_hwtcl" value="g3_coeff_2_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_2_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_2_nxtber_less_hwtcl" value="g3_coeff_2_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_2_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_2_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_3_sel_hwtcl" value="preset_3" />
-- Retrieval info: 	<generic name="gen3_coeff_3_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_3_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_3_nxtber_more_hwtcl" value="g3_coeff_3_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_3_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_3_nxtber_less_hwtcl" value="g3_coeff_3_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_3_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_3_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_4_sel_hwtcl" value="preset_4" />
-- Retrieval info: 	<generic name="gen3_coeff_4_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_4_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_4_nxtber_more_hwtcl" value="g3_coeff_4_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_4_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_4_nxtber_less_hwtcl" value="g3_coeff_4_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_4_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_4_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_5_sel_hwtcl" value="preset_5" />
-- Retrieval info: 	<generic name="gen3_coeff_5_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_5_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_5_nxtber_more_hwtcl" value="g3_coeff_5_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_5_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_5_nxtber_less_hwtcl" value="g3_coeff_5_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_5_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_5_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_6_sel_hwtcl" value="preset_6" />
-- Retrieval info: 	<generic name="gen3_coeff_6_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_6_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_6_nxtber_more_hwtcl" value="g3_coeff_6_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_6_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_6_nxtber_less_hwtcl" value="g3_coeff_6_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_6_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_6_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_7_sel_hwtcl" value="preset_7" />
-- Retrieval info: 	<generic name="gen3_coeff_7_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_7_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_7_nxtber_more_hwtcl" value="g3_coeff_7_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_7_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_7_nxtber_less_hwtcl" value="g3_coeff_7_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_7_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_7_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_8_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_8_sel_hwtcl" value="preset_8" />
-- Retrieval info: 	<generic name="gen3_coeff_8_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_8_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_8_nxtber_more_hwtcl" value="g3_coeff_8_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_8_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_8_nxtber_less_hwtcl" value="g3_coeff_8_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_8_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_8_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_9_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_9_sel_hwtcl" value="preset_9" />
-- Retrieval info: 	<generic name="gen3_coeff_9_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_9_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_9_nxtber_more_hwtcl" value="g3_coeff_9_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_9_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_9_nxtber_less_hwtcl" value="g3_coeff_9_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_9_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_9_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_10_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_10_sel_hwtcl" value="preset_10" />
-- Retrieval info: 	<generic name="gen3_coeff_10_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_10_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_10_nxtber_more_hwtcl" value="g3_coeff_10_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_10_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_10_nxtber_less_hwtcl" value="g3_coeff_10_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_10_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_10_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_11_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_11_sel_hwtcl" value="preset_11" />
-- Retrieval info: 	<generic name="gen3_coeff_11_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_11_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_11_nxtber_more_hwtcl" value="g3_coeff_11_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_11_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_11_nxtber_less_hwtcl" value="g3_coeff_11_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_11_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_11_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_12_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_12_sel_hwtcl" value="preset_12" />
-- Retrieval info: 	<generic name="gen3_coeff_12_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_12_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_12_nxtber_more_hwtcl" value="g3_coeff_12_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_12_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_12_nxtber_less_hwtcl" value="g3_coeff_12_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_12_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_12_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_13_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_13_sel_hwtcl" value="preset_13" />
-- Retrieval info: 	<generic name="gen3_coeff_13_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_13_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_13_nxtber_more_hwtcl" value="g3_coeff_13_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_13_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_13_nxtber_less_hwtcl" value="g3_coeff_13_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_13_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_13_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_14_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_14_sel_hwtcl" value="preset_14" />
-- Retrieval info: 	<generic name="gen3_coeff_14_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_14_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_14_nxtber_more_hwtcl" value="g3_coeff_14_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_14_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_14_nxtber_less_hwtcl" value="g3_coeff_14_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_14_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_14_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_15_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_15_sel_hwtcl" value="preset_15" />
-- Retrieval info: 	<generic name="gen3_coeff_15_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_15_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_15_nxtber_more_hwtcl" value="g3_coeff_15_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_15_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_15_nxtber_less_hwtcl" value="g3_coeff_15_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_15_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_15_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_16_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_16_sel_hwtcl" value="preset_16" />
-- Retrieval info: 	<generic name="gen3_coeff_16_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_16_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_16_nxtber_more_hwtcl" value="g3_coeff_16_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_16_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_16_nxtber_less_hwtcl" value="g3_coeff_16_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_16_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_16_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_17_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_17_sel_hwtcl" value="preset_17" />
-- Retrieval info: 	<generic name="gen3_coeff_17_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_17_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_17_nxtber_more_hwtcl" value="g3_coeff_17_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_17_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_17_nxtber_less_hwtcl" value="g3_coeff_17_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_17_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_17_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_18_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_18_sel_hwtcl" value="preset_18" />
-- Retrieval info: 	<generic name="gen3_coeff_18_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_18_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_18_nxtber_more_hwtcl" value="g3_coeff_18_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_18_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_18_nxtber_less_hwtcl" value="g3_coeff_18_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_18_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_18_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_19_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_19_sel_hwtcl" value="preset_19" />
-- Retrieval info: 	<generic name="gen3_coeff_19_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_19_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_19_nxtber_more_hwtcl" value="g3_coeff_19_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_19_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_19_nxtber_less_hwtcl" value="g3_coeff_19_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_19_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_19_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_20_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_20_sel_hwtcl" value="preset_20" />
-- Retrieval info: 	<generic name="gen3_coeff_20_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_20_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_20_nxtber_more_hwtcl" value="g3_coeff_20_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_20_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_20_nxtber_less_hwtcl" value="g3_coeff_20_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_20_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_20_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_21_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_21_sel_hwtcl" value="preset_21" />
-- Retrieval info: 	<generic name="gen3_coeff_21_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_21_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_21_nxtber_more_hwtcl" value="g3_coeff_21_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_21_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_21_nxtber_less_hwtcl" value="g3_coeff_21_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_21_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_21_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_22_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_22_sel_hwtcl" value="preset_22" />
-- Retrieval info: 	<generic name="gen3_coeff_22_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_22_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_22_nxtber_more_hwtcl" value="g3_coeff_22_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_22_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_22_nxtber_less_hwtcl" value="g3_coeff_22_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_22_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_22_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_23_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_23_sel_hwtcl" value="preset_23" />
-- Retrieval info: 	<generic name="gen3_coeff_23_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_23_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_23_nxtber_more_hwtcl" value="g3_coeff_23_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_23_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_23_nxtber_less_hwtcl" value="g3_coeff_23_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_23_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_23_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_24_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_24_sel_hwtcl" value="preset_24" />
-- Retrieval info: 	<generic name="gen3_coeff_24_preset_hint_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_24_nxtber_more_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_24_nxtber_more_hwtcl" value="g3_coeff_24_nxtber_more" />
-- Retrieval info: 	<generic name="gen3_coeff_24_nxtber_less_ptr_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_24_nxtber_less_hwtcl" value="g3_coeff_24_nxtber_less" />
-- Retrieval info: 	<generic name="gen3_coeff_24_reqber_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_coeff_24_ber_meas_hwtcl" value="0" />
-- Retrieval info: 	<generic name="hwtcl_override_g3txcoef" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_8_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_9_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_10_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_preset_coeff_11_hwtcl" value="0" />
-- Retrieval info: 	<generic name="gen3_low_freq_hwtcl" value="0" />
-- Retrieval info: 	<generic name="full_swing_hwtcl" value="53" />
-- Retrieval info: 	<generic name="gen3_full_swing_hwtcl" value="35" />
-- Retrieval info: 	<generic name="change_deemphasis_hwtcl" value="0" />
-- Retrieval info: 	<generic name="use_atx_pll_hwtcl" value="0" />
-- Retrieval info: 	<generic name="low_latency_mode_hwtcl" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : pcie_SV_hard_ip.vho
-- RELATED_FILES: pcie_SV_hard_ip.vhd, altpcie_sv_hip_ast_hwtcl.v, altpcie_hip_256_pipen1b.v, altpcie_rs_serdes.v, altpcie_rs_hip.v, altera_xcvr_functions.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, alt_xcvr_resync.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, sv_xcvr_emsip_adapter.sv, sv_xcvr_pipe_native.sv, alt_xcvr_reconfig_h.sv, altpcie_reconfig_driver.sv
