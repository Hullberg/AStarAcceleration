��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸�Σ�HڂͨgT�W�1�.�gW(�CpzQx�E�.�@�6��"o�0_d�h�)��"���d��?,8mN��z�Ix1�����"�x��� <��vg�m��4mF��/4$����Ҡ�o���=��X� �����'sj��alF��H*�e���w��m��H���������`i�0�c�řԁQ���!��*{�+8E�l߿b���>!i�e���)�i�:�Hx
[[��@��д�N�6�w����}Y>}���V2�8B����23c���J�Ȇ P�,��Ig&U��WT}!�C��%�	�+�cI���ݐ��f��N�W�9�����E�ÕM������h��ż����"�gP��� D�IY���D3�G��:!�����-���n�E%u��`[���n��j�#Y7�,�m�h0���BZ��`�@u7�O4r�;:�n�N��z�H�������*Aà��Jڊ��Oh�(bW�s�T�(�%`�h�$2'n�$4��֢����6��Q!���4�񉌓O�'���@�{�Z��/g?2�-z���x�x��H�o�@t<�b��I�q��S�2F��茇�ٸ�������	������2��_�@l^{[�5OM{T�,Fa��9i񵍴��4Mz,�T�ߩ��i�em=���d�`�?�'�韞�ʖ�G@�����$ \ث�9.�xY��5Y0l�NK�j��$�9�V�9�R�����уܮR!��i!r@w)f�B:������	�F�ڑ-�u�(�T���f����\BJ��5@���x�q
$1�`��Q頡�'�H~t�e�F:��R�:l_����Qj�U�Pc�7C�-���Z��$��1x��'��0Da�Wo�rR�R_�{������t;׊�_IS�<;AB:�a�<�f�ƹc�/���Rj'�k��G����獙��<���U�ۨ�4U��_���V����3�'�_� ��F���\8Wީ�I�����P�7�o]|��b��6��
˿��L���z7�$��&V��C$Q��0�m��ƭ��`#4���E����^��7Jb�� �&gKJh��!iJ�k��U��|,y�[}���z��������5�hpѨ^�?�NQ����@[\���H;�~aJ�:�QN*hڀ�,s��sg $Y��lY:dAH�uhl�PG= � L�|��<Qm$c�D�(4�zr8G]'��f�Xt��nSyn��]����l�g--i�*�\eM9�������<ʟ�9Y��&5A8:���!��3���,��gPGײ+[a����\��������x,2�F�Jڤ�Q��#R�Փ�)��Q㛂!!M�썙R�����ΰ���\҉T��t�Z��q�;H���KL�Võ���=���=���(���� �ƞ����p�1�2����d}��O��\��ǭ�.<���&�$+,�24�ql��/~�x�4 
P��48��fڣ�"Ҝx�ۍ&0x��#5�_�n��i)� �fʝ��+3����g ��`�	:i%�_?�����H)N��⸑N� ���#�8][9wux��t�ILw�������4��M�m�r�3���Vq�)�5�t�+3$E���w�����M�%;