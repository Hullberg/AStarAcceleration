��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!��ߌn��-��,�Y#7��bd��hHOE��������X���������
?F9k���.�eܶ<Yh��Kn ���1��n�%���6!Ab�CB�E�3��l2��`���{��n���E7^�ъ��4n0k��%���	���q���K�����B�v�50��P+L��n���I�d����:��ڠ˳�uS��9����4�: ��'����(>�+�e_�Z�c>�:$��h��k�H��̲U��?䞅ܧ�P���<� ��pi�.0s@��o*oZr�ҠKa��/�B ���ɤ[�r�����*2�/�]ɭ����ueUw�P�E�sG�nٰ����p%�1e'������:,^�H�~K4�m�=��P�g-zƊ[7P�uX���X)�#m���w���<��V�<.�)d9/k��^��EP6֌0�J���n��P
�Bvz'ϭB�i0�3�Je���۝���t{!0�4���gjK�[b>��������G�� ���yc����C��S���|I�(I�;.��+�Q�U�]	ָ_4���6C�I��?��8�.;�}��'%Oho�>���P`e�H�!!@�g���~����ș��O����vd�Dl�]cw� 	cւ��[�sC3��A�	*��j�t�0���0�����t����J�?SG@s� ;�A��M�e g9�?���Tl�LH�؛�S(�G\�Q6/0��C�UL���Z[������<�Ɔ���x����՜%΁���dR�B�f��!_�n�>��GB}3D�sD`�J6�fn����pB��� �M�y` @J2|��Sa��h�*����}����]C<�E�WT��:�4p�O��B�@��
�X������A�a�w�B�����k6��$���/�Y,�H�"�dv��]��js�Տk��c�.��`��zn����a���GiX�M����^���Mɉ���z�>V���7
.o���]C'3��:��b\��Qt~�_�� ߑ�9��^&����x^�:�E�Z-Dc��A��Z����+uW.hK{��+OT��
f������k�
�� Ug���'읂d^x�n�������hHz%_���?����%�I��b.���#����zp��˓�s+쎹���y��=.9��ӈu(�:����Q�y���8��UoQ��,t����W�I�z]]nA\0��7z\A;.�uwD���.�����@Վ�,�s���ƽ��P�O�ߩ��t�X�� Hu?q��JV)i'�����7(wtJ�*v�
ݕc�Z�n��v�*"'�\]ݺA �`�1�[\	�ɍ�E���{!���9=_�xpO��S�sdeQ�۸�h�f\�͌T�f�|��>0������ecL�\z7���e��4G�SFIi�о�Z�ͩ~qid~�q��T���SZVS@�E�o��8	/�1�O}O��i�B�!Ы�lKY����ߙ4�N�9������L���uI&�,Qij Âܠu�o3���� F��/�7{՛�<p�+�$��U�;	���k_i��M����Q�e�����^�J�!��H�¼��jj;��r�A qR�U{�</�ݮ��Ʃ�\�Ka��v�︸��,K�_,b|���=�P&�0��i��08k���V�>�KY��Y����h{��8�6�ʓ���Y��Ly�tE����6�ȓ�4�ʪ!'vx�d};�E-����Xy�;C+��r|���=/6��h�]�x��6U�O_c¸�J�8���0�~��� ��������t
N*��������R87`�S������V�Y��&�c��U�tkkk��,���8e���k���8�5)
��2���w$[f�h̰��񑳜���Q£y� kQ������T
"o6*�*-!W<�=~�gK֑y�	�3�"��%?f2T39�H�g%4�ȗ�9	��}).��:4nBE���+^hk�.e���&��W��bC�ӌ�n1P��j��sl-�u�~f�$>!.C�>�YV��qtq��J�85�t�IVnۡ�˒���k� ��N��Ǧf�!ۂA0�����Dą��_A��t@G���_�-��>?M~ζ�1)fpr䡤���E��`��r�--��Tl�<��8��㾟ݪD&�����(��)���r;��tjS�@�(*??5��!���ʳ�_е�Ӻ�,¼��p+i+�Dt���sj�%�����PUդ��cct g�-*�7g���bK�}	�Go���rK��х�<��6�ㄕԡ�L��ׂ��k�r�\L��@�Eϣ���=\���΄D0�V����X�-���y���bV2E�-m�v�-�oۤH~a@�,6��	B���AcFi�(��wt����^����SV�niSV��D��u ���I��!���xʑ3㏖ʅ-�����괯y�6I�X���@Al�$E�!͂2��6/�}U6aLQ��� ��7U�G����Z��f���~�2y�t�{�{�Ba8��D�ͩ�h��Pgw�9qc����H>p�#�HT�d+��?N�<�qs��Ӊ�sD��<Zf���>vrqF>���4�·-�,��uO�H����߅����� ��}�����M!�M�����3�i���d�RH�7!��M���i��BY�o��f���W�@��6�P�d�I��$�(�����^3�ΤŵЊ�T0�5���H��.�v 5�O�$?��/B��``�)}��| ����զ�!�����h��h?ye�Z�FY�������U�>�2K�-��_�[o'��j5�Rw�V4�w�#�߰����.�o
K7h����!on����ip��ۃI,qhb$�L����q:�[6����q�$��K�}�$F�U�#�+��j�B-��ZВui��=C8���e�T1�%#��S��f�9;�8�=Y2k�
6nR!�v�L����@�$o�m�U2��4zŴ�<٣*a71i��۩��)�$5�����*�M��i�	q�����@�̀������rR�>�c���3�&ngd�l�˔��w�y*���eX��\sX�$qRF^���j��Ӄ",Zt /�������_�_�r-�:�+��շD`E�1�<TJ�e�$�g���[��K����a@��f���6�BY�kQ8M�-T4�1�Wʡ%�� d��P���=�,��}� �K&�*#J�̸e�l��4�kL�q��]��6Ç��G��W�6��ֳ�c�Ӛck-��7�4$|ln���'����>��2�yD��3[)���Q+NѸ��J��gn����gc�-���ߑR ܡ�U�[���J �����VF̳���jٳb��U��ny�ugR��{]B妚�%��Q�?��6���ZH�E��*�����M1ׁ0ݼ��
�����ޤlRWZ��IH���D��!adp�_c�p_��j�}�9>+S���F,=%6,2�p���ӆAј�O�R�$��`t��'�<��Y���t3B�	�?-�O|<#�f�بL��Y,��`��)J�r)��PH�E�!����Zd}7��n+��|�����&1��� }p����;�Q=�-����`F �Զ���U�R���*�g���πV����+�M�;�-�R�d���;��٭̸��;P<��MO�����0�+�ug6����qz�龼�֐[�V6�y*�y��X��I�y9KT�v1O��Ǻ�����MsUP<�m�3�������?my������/�bms<ez�2�&c"����,A�*!-�P=��a�Ei�/�z��_Ƶ�3r>���2EΚ>7���5+�d���/�p��HD=ې�Q� ɣmiGÇ[r��ݳ�3r���ֿ��3��9Ln���{ ��F��o[�a+.N{�Cg�A�*�$a�X�?�&Lb�a�t:]�������yf!�Aj����@:(͡j�JӰ�P v�}C7p/�~�:�Fj*��X��.���Th�e;���sZ
�kwW��A��؄м��6��.��W&�M��3�(NV��]���a�c�v)I|vn����Nz�:N�+�^���"�f���o��U<�
�K=������c.;[
������:���a���
�5`��Ȝ�Z���d�X[��{Ҟ���5�#�sA��YpP<���g��g�~��n�$�0|�r��yj�f����wQ��y�,�)P�W��*~��L�@k�0@vz"f�΄ҏ�	?���_HLS5��<�Bu��h�}��rC���=�Em�^�Ŗ'9��� �A]���I�	���n@�>V�?舴�;��)�]�j��=M�W~�d��	#���8�M�I4mO�M�U�;�������n�$�jgv�a���#�sy���%De��j���tA���^1uǓ��,@*�)`�E:��3�D[Etͪ.]���� +�Y�>t����:�qt}����IOOPs��*�Hy�W'O^�����=�_��ʋE�՗��,+�&x�����bH�7ދ��cg"��QƜl�RR�CQi�L%H�0L��p�ms��ǭ���m�'=�&���$���������?� ��Q�/���Y��k�(��d����'���m뒂QГ����Y�=��G�#�=��?��vSs3^���a~�혠���=�y� ��F�D>%ʈ���-p1p��.��.l�YWIt��F'�y$��HF|����������SK������$e�cZub$v;/����O0���,��"+{;��X8;Dy�P���
��!�
��ﻬi�f�*�^8�K	��N��18�مf%��?*��y��~��&/g�孊` ��ZJ/t����,@��%�Ʃ��WUG#,? ���d�b�����x.�qX���6�ED��Z971�~�ivՌ�wP�p�ts��m2���}��� 5x��D�pZ��r�p?+0W��E�.w }3 ���z�Z�{���}�G��dd����o�v��a*�7�� h��a9וA��K{bc7��#�Tp2��TF���,ǃs�*�_R��{�W�T�TY�Ce�U�=am*��gֿ��ﲩeW3��gn���ϓ�j����E�ĽL������F�|��;���}^� �`�<(U]���\��1c�U�oY��/`�J�0"|�]F=b*ۗ�5�A�.�"�~���f���i^G�l��+�����qE�*.>�ۢ�Hߞ�8Z9A7x�
���������\��#��Q�O��#+"��؁�!6�ct�5�Y 帲*=�`��;V�ǈ�YM$�y�`z��E�O5����u���AN�69a�l�a�����b�,��e�U:~����������{�U�h��
�h��
�?螔��s�|�v��Ύ'�,�*n���>ln�'��E	*��&���>̤#�pZ�ͦ-���O���y�Q��s�5n�_���<��P�-�
��.�S��]`�9�"��~%��/޻��F�x����A�� �) �׌�� Ă�je�>Ɍ�����KR-F9�]�"�cmJ��}(�s��f�#��I~w�U�������j��i��!
�ø:����Fj��*����:⿬���nz&_�}!K&X���Tz/z/��{	���%\&lR����S�7���`�����%���E$*"��R��XIƑyc�4{յ���r��n�4�f�9�O<�_�X�)�y��"���;����"��}ɽ�Ѳi�Ψ�����Md%�[NW�%hg�(�1�,W$��ʣ�Cm6�s���?'��xa�WMJ�Sq���G���-w~�d�.cK�.�1�"�-h<�$���_�!F�����8�9���Qq7�.s>��n��&,pK����1�7
��64���S�]H`�~\�V4H��cƶ��=r����1�t*����
`pXCvU8�?�{��.��;y�	_��04�Ga2�eD���ƪ����`{e��x�>DER��<�/I�5q��	�4�"H,����E��e��
��~YJ�ooU��-u~�u�M�������k��AtKj���ئx�NP������?�
^q��3wßĜu	���"rc� �4Nb�Ɉ^vº�����F/��2��R���(/ǔ� K�x�Wl�c��qSt�Z��u�{>��J֚7Q�P����@�R� z�=F_�����d_;Z=2�<;4j���{�?@�C]=�e�X!y����,[T�Wf?Dcm�W���VLIS�+�O[�zp� ɼ�PGh0��4!�w�`����?�E�^`�`��@榕ê]o����GR�<��yr��;�J�-���ĹD��;5{d� �JY��31����0:񛟂�l��
9�a9���B����^�s(�ۣ�LnX83��}m�yI|N�(&��j3ų�ڤ���2m_K���,[=�qX;�>\R�6�3j.���FTs�G6����8vI�[i��Q�^?eu`�)/�ya�r\�����jh]�����ʿb���E���Q����$00�䇴�c-!��?L��m���2B��d�!��жt���ah�����f��(�͸�+F�xE��A�����V��T�$G�2s��G���-a�r�\��m��5�	�	�:6^�f뿙}E�rQ��p]��K*0��V��;�n��j�.ꒂ$�xW!��
4�%�X��̇���Z��YƖ��ؕ#h��/�9�䋎Κ��w"��	"Į�Rp>�C��vn�����	���n�8r�ֻNT��`3Nu��{D������t�o�K�1V�7=P�0?í~�1��*R�\���\����N7ީ��8lQ�X�T�9]!}�C�
����e�ۺr+�e��/��D\��g�6�]��_�x��8��N%H/��.^��M�����4�5����R��^�pG�(]���8ԁ��/	�@��C7�ڢQ@c��51ݓӏ�.eS���W����4/��z�GJ,���h%�s�Jg��M%�c3�<��w�+����r>j�;�0�EYa�A'�{�����M@I��'��6�t�_܉�ϙh�- ��:q۹��M+�G!�{g"TR���S�q8D#���dl<Ý��g��6	�.������̙vݑ����b�(F���<�Nɣv�
gʑ��C�&^��o�>��2|c= �d�Y$#kW������RS1�&W\ˀ��89�tN�o1�ؠ��~�b��90r�
x��"A&B^2T�Í	%s$:��_z.�zήP�e'�q/&j��������l����!eM��[еsU�Ҕr�~����ټD���?h.ݩh^�����\]C�&8��^�X%�]y�$��cC���N#���9����X�Jc�0ՙxh9�� ��e���8㩳B�	q6c5@�L���2ֵg�%Ӷ0#�v-���8��
�Fs[�D �]3n�C9������Hs�R�ƴԍo`�ܩ�X���%u+�b�?�:u^�E�P�ub+�^4�����ұ�֢#l	��k?�e��+�yD�� ��;�Da����f��p�X�M��q�����B�RK��(�&\���	+T�6e���V��ɽEغ�p�� ���!g��;c_�ő�0\6 o(k�<�Ʒ�j>/�0hD�~ZVxךix��o�5��O����v2�t��M�/�ؼ��ϯ�n��	�g�?H��>����+Ns��nJ{f���B�L#��8���U4(A[�1�I��Ύv8_�o�)�D��\֞��T����i�����D�[%:����m�2�~,_s���+f"q��Ģ��d�eFʚ_#�2��I/I\��vdY�4`딠�D�v�ɭ��)���ņPur���[ ���֬B&
f�:��d`7Y��Ofz1�}%�:S;�$�v�)t�<����I��sj�n� �r�z�@.l�WT�q��~����i��ĺRs��[�G�E���!x����L '~g�Ǭ0��h�XfG"�(��c�q���	�Aws�	~YQ�ō��EP�7MH�	�g���p����#DJ�w�/;)(���sY�P؝U�1y:�1��v_�@-�Q��/}�֜��ϔ �B��)��D���K�_�,�{w���]ϖ+��n�+�T��//����=g���?g����=�Tᱨ���A��ۍ�h�����nP�3�5�}��<@S��:��W��ҝ���;cs�2	i��|w./@q=�4�p�L���J�$ޯ��k6�xv�����*9l/8_�?�ҟ+9�SQ�cAa�_����ՙ)����[��� ��\���nmׁ�(�I�#F/�=��\q�㷢4^H�S �e�Zx꾴$�bA�1�X6��Q�ݾFtL���E:�����_���U��j�P%��7���\'��������!�Tc���L�@}��b5�r�DY�K�o�2�]�|W�'�_O�����PS|:��~��L�(�y���[=����V�	�dҵl�k�_J�|��뫅F\�-)>\K�Ҹ�ɱ޻B z�\���}��9�#	��<u��X�2��0�h4:g��� 0�D�J���w���̶ںNrJ�P/�}��m�Sy�����A�<��M:݊9(%�^���P�n��2H��l�=�Bk�
�u�I�u��Ni�,�l?�z;���2M*C��x*�z(�N��c��movRbuo�j^&W�լ0�o����lˡ1���G�olAn~1��:�v	b�S	I��4M�Pzld�R~��M�/���:����4b��j��	kj-mn�l��
	����ӎN�8~���41e?��Ƭ ��==l��,�X�ęH`ҺE[���c�/����M�|����@B�ֽ%�d{:�}�����]7���TR�ʕ�4Fm�`Ty���8"�to5����VX�
�1�'���j/|%�d���l3!ͯ�X�,�Md(��#�t�.���������v9cg�Nr,AZ�����O���h!��**EC�~7^3��������w�}�y|կ�\���7&'\-&����(�5;���c�<���������bF&�îqU���Q��I�#߷22N!�PL���#�!q펇�;r�Ҋ���l^G֎�� ��.�20&;n�Xz�*�p%`�*m�fG���*�W����"�u�՘0�h4��"���HA��GC{)�ŖS�c�/�Tz;Dw~�3�TU%�ʆx�cp�Y&|o��ũ����Wټ�Uy�C"E�S�P^9�� o=��Xu�> m~�1~�es0-�P�p^��p{�[y����OC�lַB �]r�D�޽ћ!AՖKYEl�߶��-�֌�ѹWЬEUc�}�o����H-�*f3�R���T�KX�ѹLj ���"��U~��łN[q{���g˅�+���Ut����?T��������h�|�Ѕ�l��N�&=�/��,}��G@�'�7��ˆ�#�'n�祿>-d[$�2}$����[�%�������x�>�9E^�ɉ���-�/uq}���:�K����^ɉP?h���q��i�*0��<���G��ж������__V�Cy���5��>}����C�tA��<��iHm�����P�� LӜ�H@
���`ǩ�T5T$�/pj� N�]��0/>���%d`�m�����ЌI0}��.�&��0�)�63�����(������!i���#�{#wi. �n�6q!>4,ou���W!2 �=�r;HT��7�K���gS�j��nG�͋=��/�w�rN �MZ#�?�{F�?n6�يIu"/���j��]�#&BW\����]r�6��="�dDڜB���(=��r�达\��p���W2�l+�~ �� ���kE��aq�}�N��� �)G��E���V�༔<���=��wߪ5L%���֞�
j%�㔉���ڪ�)���qt~r���2�����j���B��R8TX���F��H�- �v���B[h��+���a�q0,�d�hL�X�u6C��6���Ĭ�V1�	Rs�
��s�ʅ�Z:��X�6ƞQ(��r��l;CBo��kD���*�R?΋T��CF��e��Pve��PN���$��������T��\43�a<�:ډa������
㒤L�g�V�aBf���q2�ki��I%6��H]�8e��8��;��*ŅЈ����I��w�o�++��PC��a�u���Z����W�X�|��
�Z�����4v�s�mE4�4�:@�8��=��NwA߽�!_U�	�/�k�G�*H�s�41,w�[�Y zG��������psш׿
N��N��S3t(�c��-�ʖ�V4q+ ��3��Ä���m뱼��x���<`$j�Ꚇ�?8{r��E#Uv��O�@�-�G��)�h;1@Ñ�Ro.�E�~�! v�_�,9Ę?}5̹��:��	�a�:�u�����:u��-�TыT��'@Ǘm�6�!���a6��QC���Y�G�m���y�c��|̵�0�@�|<�Ş��o��yBn��9y�8,Tg�U է%~I�M9%�V���YV��z���`2Z���D��*밦B�mP�#�eqtz��C�S�E��'P>f��s�ƿ]�A	 %�]nF���Բ�h�9	,SdW1��v��#�!��h_��(�k�[��ރ��M��g7�I#Vy��ux����sl�?��K�(�~Q�|����Z��n�Iv}X�UA(�`��Knr��S��w<�C��	�^INt���,z�-�r㻴4$���8UQj2�9��3'8Cd����.ߵ��Bg�8�!�z{w�;�|^h�e!��	.A!K8�8�'ߊ:k�"����§E��7^#�K	�����mC'oWhE��-L|_Ӻ����^
^3��O�~�r�#�r�'h�H�ဲ(�������;���Ã�3ݝ���p9�T��&��@�Z�g]�f�^X=`�#d�2M�c$�"�%�w��[6�hz��C[��?}&~���j�D����o�t�,�M@�b;�tGv��9�k����b���Z��7�v�����)C�a����R�lZ�����]!@�U�a�7=�k�|r7*D-l�}�f�/1)#���KVF"��[p��BLn�n5Iٶ�:(Nɤ���Bn����?N�G1�E����h�����Zc��<*�(�x���s�+�&�r�$�Ma���P�δ�PL8���dW�%B��P�����	�����$h0�;���p 2ad� ?��t�r��b�@��Oy��pʋ)��/�?�\|���*'����n����V��3������IװS�Zv�z1������z8s{20l��|���l,��z@eֽ�\�2>��:�^�˨g�� �L�����60���[آ��a㹼��!�_��c|q����T
���w�YM
�e� ���e$�^;c����/�[@