��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸�Σ�HڂͨgT�W�1�.�gW(�CpzQx�E�.^F�tZ�����t�I�k+ǉ������]�+������d¬��l�y0��FwOӻ|�a%ZV��
���~z8�q��tqt~�Gq�H�Û-�H�K�lW`vp�@�h�2�Ն���\w�![�oBy0�'2�2��<��3t���T6�jeXTt,��Y�S��@�
$�Qk��-�EHg���3K@`���S��S��N�%�ͳ��M�{��;�H�����
V�P@�Y}x���0wO����?`*���|�ݎ�vn,�B>p3OoЪ?9��	��pS`�C�֭�Q����� ��rjG4V��s���:kS�$I����1{�+���(A6�K(�C����bIV"�&U�׿�� GLҎ�O[Wb@c�ބ��h�h8t��M87�&]�^k�j��u����]�S|	�% �͸�������+x)o� �:Q����v�k�ͯe@� �i#���BC|�gKH���zf�qCW��5tj3v��}$޶~��sM�ߔ�l�/�]�Q�W_��w�Ny�bĻ����ڲa͍�TgE�^�?�6=��z� Z����U50>���'!�9_�?�]�ʜ�W��z�b����2����g ���Z���U�g�Ɉ?�\�IN�z��p�[ߓ��� L��!;��u(��8�������!�8�@B�t�?r.9Q�L5Z|4��t�<q�]�SMl[Ff�<�J�Cm�3�t����ܬa��K��&'�u�|b)�[��x5���<��r�l���,�Q�P�w�""A�S^s��k�.��] E�#�����~.��f�8���|R���c�g���
`5�A �= �'����^�A�ߠ��+���T��V�1 /�����k�%[A�Ou̍�#��T�~�T�R�#��`��cW�1U��~S��UA�*Н�XW�\Hd�V�l��\��� �ԫ,�к�
'I��jiM�\i'���X��!�M�5~br-�0 ȢCМ���f��r²�uըE�vV�z��<�N��B���ه���
��ܢpl��{�x��j����v�r��"��x�J�i� �ˮ�F���&#���Z:�����#V��s����m�&{	|�׃���k�Q��-�-q�Z��,O�μ=���_Ѵ�c���6MS鸵�L5��v]�����W���|P���%Ss��dq�߀f.ѱ���BNyJJ*5�oa�t�n$�����7�sU�Y$�����Ե�ύ��b4�'a��6	R���O�e��҆O���g�C�f���^B'or��l��`Y�{��L��_2J��r73�ݭBY��AY�a#:sLOH��O�H(�٣A�`�X�XH=s�l���m]C�����"��c��i�ӣS4�0>]��\�����Y�N�.VL���i�<g�
M�}���-�d ��H�����I&�i��0j�ϔ�Q��6A{9�<����.]���:��^��;���Zhȇû �࿓���9���ɝ\�ǭ��z�{� S~����=�ů�b `Vs�q"�L��f"���Q߱��e�~�������3�fPQ�9���83�����+k'�)|���7�_�7���}��b���z��	��&�o�x��-��i�1�	�<�5b@ü�8���W��?�`��W|G�~��Oҋ�#�`"s�ϣ��j�����s����Aa7;%��Iٹ�e�OjN�42�B��DP�i�wٙw}/�]��͚����