��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!���ff�a������b�PG����<RS�%�9�k��M[���:�tV���8���Ƴʍl�� ]��N{w���Œ�C��Ȳ�Ѣ!���Rѷ�!�#�� � Dn�7��(3�S/-ifa��$���_K�,����Wqrzs�>h`Tg�~��Ul!Z����ȿ�9T�=y�׼�*��9v=���	�t���<\��}�R,�!���i_��>�*e&t��R^Ĥ?_�^���P�,@���\o�����n~���b�i���U�������j�����%$ez�vst�y7S��z���BIÜ��4r\��h�jE��j��� �J��Yf�Z:8k���z���(|�V&w�J�� ��`�A��s?��x���}�<�y�Tr 49,���N�e�W)-^́�S���k2y`�d��Tw�N�S���k��>�HY��X��)��y��e�����,�6H�;�|��Sшl��H[i�:�^۸��{�"<\X��M`=��T�7Y䅒�d���� ������Q�%��Ɖ�p��<@�<�O �5Gk���������}�U��8}Ǐ�����u蘔�2(��Ab�r�9�c����
�R�P��fG�(��֩6��Y���64��Na�ߢ���	���h�d��������JK����RE��8���G޲N��TAV�ؿU�7$̺�^î��d�Am�x�z��\�u��u��P4>��X/�Uw�w�ޗ/��;VN�2�^�.�Xˍk���<���[�o:�i����QK&O�l�8�.3�����S���Ѩ�X����AL< d�����L>���S1ë��Fs-G��D���u+�c�M��$��XøZL�>�}���Gh���1���� �����9n����*d��HV��7}oy�+�jgn�c��`lwvЍ"lj;6�X��Zs��ҚNW��6h�?�8���$#"�����7 �k�X-̦���(��kT�"�oQ�y�>Mw^��;��Xș�	��E-��ޏbH5ib	U�d/�y�䗼��x�����r!W��:~���B9+����"�N��#eCA�6?/z�g�y�g�8��e2\X�rP�BZ��1<���qn4�Rj��=���q#���c�.���bܶg#�h%S��\�
3S�
G�8a�����3�_'�Ii���2]A
Bd�6ør+�����	V\J}�0��N�G������]���m*���rQD��Gy!�˶O�U_[�Q�c��׀��<!������[�����}]��YO���b��)T�zHDO.r2\�?��1-�^���σ�j@6.Z�p��Tzi�.�č�T�.E�-��-�`&IhL� Ӓg��}-���1����*��)�ԙR�[�g$=���So\^3&�r~�\��uv�Ȳ�AN����<�������*��oZ��K6ԓ��
��;��E�����J�p\ZF=Sc5�*۪��Ԙ+<�(�S-��B[o<~Ҝ� ����DpC����'t`N|��I���^�nP�]����k�"%���zg��sr��݈]N态5�&抇�5̥�lv���](]� ��wƟ<+aGۘ�#�e	FДz7�Ơ�TZ�J�w���hz���o-�r*D5�qЬdpr�����?l�`����W�Ju}vc����[����_��3b+�?�2h���\���>��4�0d�N�Z{G�'�`M������\<z���w���J���p|���ҧ�}��)�,��y��G��!m��cQ~�7���k,d\0y����+��U!٘��5r��y�q*��o�9�-�u�V\d��K��f��'�[4�\��a��7)�˝�X��3e��v�>��+Ϛ������@���~�z*����2�r Z#�/��CK�Q������]�`��	��]3a��g��Y(Hx��ӌ�4��!�!��r��7U��R��Vӄ}7Gk6c��,���>�7P@��1�hP��z?FЊ���]�̏׷��G�߹�($gs�+*.�1���>ڇ� ��:����޿l�����bU����Q��bZ'����z�1h��I?;�0nr���SI��I%��U�+۞�(�B�����[~�����-{��/��&O̻X.m�9ꪀn��'�&E�B�K��|�>�10~�Q��gãs�_��p��X�^��{���t�w%C 
�)������*_���BŹ��5F���<���_;�a!�f��1��5�U=�,�E���&�Wr��)����,�[9�K���x�;�Phvt`_AsYr� ���J�cD�{fW=yݿ�l�enB��y#]�������u��i�נ2<@`�w�oOw�Ŗ�6�LV���HK�X?R�'�Iq�|E�h����(6R�B��E{!�����	��P���yڿˈb��l��͛c�ǱUJ�>�KE�Zn$�u�M�?:|����(��2|��t��6��(4a6�9�����h���0~`�<�Ȗ
c��(��L��"��ͩ��rR�9[4o�~]��:��9c�$�N�I�?f�#.ƹ��W��~�-h�/ ݛ��O�C�Lu<�Q�v~}�8��*�B �]|�p�?'Ե�ơ4��T��7���Phul7sɝtsY`��F<�
@��uZ��-;b�"1\p�Q��I��6T\��+��r(l�Z�,,�D�^u�T(̼�r�5�?7���b�y},�hQ��r�K�~ɇ-Υ�w���s�_��t]���ϥ�l���Nl��9^h���6=��Z�Ui̛�\�PX�|��4 �[S�LI8�+J���))��E+��I�Z�f��Ê/���m���S�l�\Z�, &>�ͷ��c���$�[��,�0�a���i��u��2g�	^�㵧��Aa�sV����ࢹL@Y�.z_�`�,�o�6I�+�(ד\d$�Z+v���T8�:��-�g^�Vmt9W��vP����J�AW�W?	X�s��7It-��	t+i��*N��,��"%�[�Q�1�Xp�����M���&n�V�Y=f���}Nb�}'	C�@^�@�����lt�-�������%�w��h��MJ�%��2X���P�Ŵ�9�-=��e��F��$=/E`�����?D����/�p���$֕ɩ%�g�oG1������fc��2���3������_Dc4>��U�7&ѩ�ɟ�>ٸ��`��{�r��������z ��)7�}Oi���P~���~�d��!Љ1nV* �d~�(�t-1"���`3���S~qB3�/���m����T�t[5h���X���G��ՄMx�Ѣw(����6W����GRhN�&�P��0IW�� #�h�9/K��-��ǂ!�G�E[���>�&5���9�7U�$�Q\7䢯x�b�Ԉ�ϕ��w/ �?��-zE[�!Z�m1�i�&j�SK�C�/���
iw��@���U6W�PU0cj.�ѡ��Cd��l�7�b" ^n���P�7Lo�+��?�]ݷ �H;}A�
cX�R95lQ�Ʃ/y"�us$*)�nO�.�bgNጱ��Z���iE��$�.�P�a�u��G*�:�,��4%Y�UN�`+4A���lB����G:���߾X1�G|G�ښ������Us_���j�ݭ��I�[�ы�j�읏]���v�2�r3�_8��CEc��ڨ���3�K���/�9i2r��=N�{�����v ��=a]}�8Ͱ#nHp^jڣ��O�D�% �a�G?�y�����;�q�TK��h��6a}F��B�z�ބ���}	�5���D����� ���YlH�"�1��.�:�;��[*m�ƻ�Q:='v4�A 'Α���+�0�s�����:�{�+��5��%�C���*	H��r�	���>�u���}3%@����[�a������)���	���a��r�K�k4�J�e�F8Y�(�!b� +��_�G�	�(�X`�'���h�D�����������MӫT�>?����T�1w ]̇wD�C���oP��3i��aI�bCZ���5�Fǃ\ˏ��R�
*s ��P��΅�+�:�z	��%;.{f��,���g�M�ɋ�2H�<eo������먡c"����n�=�:��BO$T���]���M���ɤ1�xY������6��e��C%�o	�O����lrS|4E���sl˹�In��z�-q�L?�d�E: �H�c�x��y/D�/9m�@���Q\g�ڜ�>��K lS�sv�0$�v"�H¶c��0�Ӗɥ�m�E�`��L"2�Zl&� �J?E���w�����z���VVfT���������_�sd$?�kg�L&�k����(%��"B�$�ݽ���e��1$g�(09�������#.�ǭ'P�»ؕ�M�|�u4#S8�y�3�a�e�#��rY3����S�{�mړ�+�p���/�Rz���N�}�i�<����n�:�]	j�Z\�f���Tڊ����0NF	]@.k��:�=�9�J������������<��8���b=Y,���Uif��kfs���� b�,��a�%p���un�'i�;$R�]�f�ɚ/G1vC>g�����K��0|/<o ��RL9��iDp6�Us��cR�������3	5i��͏�>��MR��?��G���h>��`U?Tkb�RY?�w�2�M��Ƀwdn�yp�O�qCqz=����#&������߿���ޟ�'q��^�i�mf��j���W-�1��"p|���N^��jR�Ù��/�f���g�F�xr������(����?�P�jXh!E���?;P�L9���� �R(�D�������gaEl��H`0�óǳQ`�[�j�s���	R�%�v[U+c�O���>R0a@�;6��i�Jژ�ͮ���ˉ8���oS��E�,�Y40�ϡ➶��Rg��U��ў{�\3q���ea�~PMK�7yb����I���ϡ���͒�ߕ�R���֯LB�O�@��uV�����yO�
X�aOEU"��g�5����^��-h��0���RE�֢CtKE�����сjbur��|&"OЎ�)L�4�i���1�Fؔ]�/�(.�!�Ƒk�/=��|E�� b�g�'t�����Bp�+���/�u�.�ڡFX��+A�����M;���%�﫻���jn��-qS��4VG7��/��hG���lc�aw�V��,��wf�M����n�������۱L�M�R{��K�ѹ��C<ۢ���[r�?�&+_)����V�n �3�]Y�.���
`���Ș�[���3\?v#ڂ}�ré��{����qI���4E�m�����U�����чg���(�k� {��
..)N�pÍ�۰27K���e/62&7��%l�3)l2\xYE����,��p�;D�,f[��CB~�����,���3qvBB���C!w��P#x���F�=Wc�*�I�]�Ʊ���3Z ]�~�3��K@4�
����UH�x2���]����n�NI�����
���y�P�6��;U����D�K�����C1�I>�f�����R�*r�.�B̍x	�.hd�G��O��R�f�6�u[�7*#T�.�y�Ƴ�EY����ڀo�v9q���tA�D����q�]�?پ���ōD��k�V[��\lfq�]A�*P��G5�Y(��y��X~�.t?�1�z~�3jV�±�F����%�u����#�3�f(�,���s6�:B��EĞ�`���j(s_�u�n�ؒY�H�7�c�#s�~��ܶ�V��yɽ�t�%�Y�/�7�Ie��t��l���FO���X!�pOqNr3�<Ԑm�\�T~��5S���aѥT�5%�# ?��>1���J��d�ys�2���:��0ʥ *���q�1{��>�p6�����U������d8YQ'�w���i��
�)6��Il����d(�-"1��O�u^^^��˟�C��)�K~e��Q�͒䦙��D-�����+^�2>0�ӗQNS�^�Z)���yP3��^O��jg�g�,ӏ{Atp� q����o�n��}�g*R4N�<����
���$]	J�K��d+i��p�M8�v.�ٓ������ñ�/�/X�BE��n�V0Ȏkec PEc|/m0c�.`��I���W&��^�Ft���Q{A�q�ͷ�:n�6�*CQ���O�q1�k~uP�[�JBE��.wd.�J٭#�|��'@��[%�C �븡�u]��7��:!���=��6���U�a��ʏ�ss�q���-7��B�IM5����z	����&cx�G���� !��=�Sd�!�/г<��-b�	:J���_����e�tw��>�saF��<|}�sn�y�W!�=giuU�r7q�����r���\��ƈ�>�֬U�| 끭^�P�[��g:[����;P��t��r&'`8)I&w�&�F��,75�
�"�V�p��0��^-����צ���IM{���jbj'�I�`� JJ�n�CL�ZH�~��[K2%bq'Bg��ي*����^��+3q��&8��w�m���9���,g{�d�`�D#޽Cy,Oc�8J�H4/q��BK��I�^��V�s99.�}{j5�;�.�l-l��0�>�s����V)O���ۭ�̚�}k��Q��ӯ~I�H�X���å:�u��I�j�}݉�A��A��y�Ԁ����~Q a������^������4ž�;:r)��*]�������ܦ˅�>~��Ұ˼5s�a��}c������H��2
|rf�U���8GÄxyY���L^9&Y� At�]%R*��r��Yz{��m۫ն:���].YWak��]L�L\WX<<s���@��Eʥ��ciuҧ[�i�T��q�6��^���uR��I�"�	w˟js͖��W��#G�(#��Lu�� �y��%9z+1>���V��K:��_="��?��np�E3O*�C��=t�p��P+�.jw�"t���4;�D�� @��(FO�vLE������J:T�**�$��X�A�ׁ�w��ޟIu;���"E�0%��������S��֔���(�{��3[�<D@����T�m�a��8%���T� J�d�÷���!�Yѵ��3�!�`��|L�F�ih�pSCZ���J�]���`������Up("X�T߸�ݾSA�����@�H�g�(��8�h�<I~|z�7��e��#1g9��0�5G΄O�K}a�AG]j���e�ܡ=y�	����4m���TW�)���q�(��;rǽh��e�.�"����+k�#�F,����?����W��l�]Jn�J�����u84�&�nf��N���m�ӮjE/)�GB  ���j��OoXQ-d�i���f�Pe.�f&_�u=H�~��+[��\Tb�Q��9��tѫ�`�iV�+��>mOO�*"Bܙn����8�?4X�$~����XLcg5ď~	���	l��vL<)�k<��� �-]�Tlr�@Ant����d@A9���F���)4������f��,е�N��N#����u�Q�񧘇I2_	1�4����� ����^Krɚ�{F�� �ZN�%.-nؐ�0� r�3�'#���k��3l��T���8=�|��֓4�LWBy�2�<3D,��b�Z�=�<E�s+U#�����/F�ɩ� 7?�k���M�,�?+�11J��iE�A㙨xf��r��L�kB�5�P5�&��:Aй�&8얔^Ň+���?3��z)�s�Y�۝u���'���"��������$�`��������9	�L@���E�c>5] �=�Y�I,��b֫��Rxu�[���CW� ��a.l���q�����~_QM���v�9�x��*t��NH�g&TK�=�y�#���WE�v�����fq0#C��Z��g��[#�J6NU=q����BC���28��\���%�G��K���!İJ@X��1&9
}y
Z~�"���H$�����گ����F�0e}��.��Q��=�}�ٗ��U�5+A3:������Fxْ.L���A�O���؆��^V�w�9/BU�U�P���iMm\d4A�K�w�����/��7���<Rڋ��ZI��Ά������1쨠���
�T."��:((J�O4(
g2���S�I$�ȕS��i��s ������jS*�շ�G6�!�ZUvJ:T2 eh��8����!p��D�/��Y4�gxfj1�UǢ�q�1�|��*�!IT���ք	_~�����M��$a�dwkKx���+c}4-�G��M^,������Z��4�>�N��}�WH�~	@�2����<�͢�p�\��d����5�(�kmy��u�}�I+��K���*]&�~/�RHpQ�zX�x�{�=/o�g�Ql�-G��-bnocu�;Ӹh�����L���?�1���W�7����S��:�W!��ӻa>/{2���?����y(������5�>�:��ކn~3z��ΩF����x��\1�Ó�VŔ���A˿��7�~�u�Eu�{k�S�����@j��c81VG�Cs�w�Κ�z �-��06_���{��z׽�%L��Ƥ�e�|fh0m��$"�:�|wM�y/S�uTA�<�ژ�IC�~��r:�y���feBa�jãs�cHD�^Q5��W�e��b��Ub7�)��DzńKsP���{:I ¹�	z��g�:�D�����	��K�\enF�t)�����������~��=���!x�mW�5!R��\P2��_�(9\�dD�Ȑ�� X"�<u��aQo��%*��G�j�5���Ёt��H��@�hPz�]�a+-xk�9��Is;�m$�g�E�M��_�=�i�ƕ��G�`�Uf�]�5�d�ч�"��S�[䷻��{����m�k