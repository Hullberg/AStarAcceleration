��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!���d֏�q"ed�1�kȞ1�������@������]f�Ȩ��fa0{T>q.�b	G�(9v���ק�^!���Oc�T�|��z?~3�X�f-��������Y�D�հ?H�	3��7qo���쵭yp��Q���:2:W��(�LH�v�"GL�,�q�U�/W�4�ԏ�Б���# �> ��3��������_�i��}�v��+)>�e����bkyޤc�M/E��U����c��[�)	��΢L>��^	kTʥp|��.*��wz־�,=$#�c�P��6�|jGjWi���D�5�*����h�v���]�&�&��+#[�ۓN��@������rW�μ��vׅz��=A����-&$T��hElYXp��4U�p�֕��=0�-��W�H�5����I&1�mF�c,�C�Z�U?jX&��o��4��}
Ip��nA�N�d-dًU���Q9�$�N�2XL��5Ғ�����|�3�H�)�����y���_r`�i]�2��%��RL�%F�CA����5�1����R_������� �&�E���u�]�s��J�����J��7��S��;l��T�t��8~��Ầ WK��j�^�r�����KVy��}�ơ�E��%Q��ͥ���<�.�����/����K�a �%2�i/b���n�oۖr���AY?�0~�'��x2����B�ӽK�f\r����q�Y��;�k��ç�M��U��ʩ�6�t�܀�C�ܮ���*n��,&²*�Ƭ0�6���p1��ϟ&(��9
l�Ls:.�u���Z��D*�����%
h�	J \��֊s�1o��X<b�f�om���6�<���=a�T�R��vA�̇o�-?�M�l�~?Ys,p��S3n�_�������3�Q,�^��e��$������S����P9�w}�@��H/3'ad�(L��:�cy��y?�՘\[2���:�����V+��h��M�����I�)�u$ֹ�u<�:.� �ř�E!���E�̖����c�z+.�N���/�^���2�����3�̖��.�O�[��L!GCe�\�(>q���qS��}�z\NT�s��J���Gr��Z[]J�io��� �>0b�uj��4���}:O�eW)m�����_'��v��yn�>�w.�7a�l{�ܬ^��h����[���8���"�K����yԡ#��[��"��i,��P�r��"
�؂��hM�[ 'C�(�r��Ȅi|=Ke�ޛ�`�6��3/��_I(E������&q��v����ɚ�|��+1'���ն�����	�C;�����EϷi��\5*�>�OgV�Ɵ971?���Ey�8���ꖎ�5}�yH�wLs�3Y��Fc @4)�HS��a��2y���Q
�tFβ#8�!�F���/�6!��0N�,�y}kQ�K�>Oa���Z� ��tA�eդ�b;�:e�AɟA�]T�f��t�D��������rƁ�8L�
�T�e�[�����?��C[[��DH����&V��j� W��V�{W���n�R�v����mg��r���܆��ض�6֠�"׉�V�h@ -�2�~c;aT�+x[�(��{ D�.���L��eUs���2G�qi>����A}��Z�d`~M�o`N�� �o!�C����18�4�Ρ��' ��� ������}�׸���'�7�詔s�\��R�M�������@��3}�r�k�͇�?2�bvl�?�N�1�a ���:��|�ɦSG�`���$bswD�8��S�1y�D����E�akI��>sq��#ۅ�lb���aO�8�	�ʹ�L6z"�0NIA��5re3`��O�m�����@.\f�(��|�iҬ�fG>�yG'q#��-��t�D`��Д6��NZ��-���F��:�P1��I�߱�V��kK�qW�Ϩc������7�~!#uJ3^�+|�3�1�?z����a�1
b��֍.��#|�9ǅ������P`�a�J|�6�5�;���@�d�H�]�v��L���'l����NS}�Y\�#a���쀧�sGw��M�n֬�Q�B2���l��7���,�
�+��"�S��G:����Jڀ�me�����&��Y�y`��Ҩ	����1����H��2���. �*71�V�(����߁�M�݇TH��Q���������Յ6�7�6�ͰʈhV&�/�����6KSK�m�$��H:Z8qŚ��G�� ?�m��O�B��m���X�j'�o�D�V�5:s�Kn��!��=�mZ1�9\}���u�y��2�9ȆfR ԓ��+A�To��?�"���u꒒��y�$�`� �u�0��E�tHAL[B�{���L�IZ�����4�fO��yQW^���r�o�Η�3�ڧ0,5�Jg��B=m�U����
@�v2`f��U��v
�]&���C%�L�X���	OqV�J g,��r'�rhtQ.մۤ�u�"� _����x<8��L%���Z�P�P�u�ቬ��A*�
��;�T~^��ѹ��V�c�x��k`�{�l%�9�� i�IUŮ'i�W&J2�>%bH`Y�����e�Ǒ��:Ri/(��3�����@�^��Z�K6'U]�5-������;��޽���{-�����ե��9�m����M�'~s𑕺�YJ�P�P��6����ٮ�A+�@Xbcfe1R%�����)#�uzhu�_�"��i#=Hl���!SΤrj�$�(Uڕ��0��KM3`��[� �]*����(��R�23�y3��Vu�_���f�4����g��j���P��L.䛃�}���iJ�a�y\J��V���k�6�Y.#f�������s�e�X�'j�P5<M%P[tϽjQp�i)��b��OEٯ��ad�m;��� 6�/ؿ�|�@?`o�e|���QY^��K�|����~�=��2��J���}�%�E�̔ﮛ�.��.��Mϔ�#d����?���qW��\�J����|Y����M�ȏ	�:�Dip@\��rÌ����H�+`ծ��7���8���Qa��ϡI�b�a�1��z���h�c�롖^���!�TJ��w�I0��Ý�{R1[�%�����8��ю]!���2��1�UJsH�pM:�$EH�F��e�`���E����2A�9����J��v ��0μ��	��6�q��PCv��KD:�tτ�}����ݵZ�J��R��5��ن8�m!q߹�
�w�nHP��ڇoe��pcu�5vv�ێ�Lz�J�F#��O��̈́�)�,+l���	� ��;.G�Zg+��+U�ş�M(y�;]��7�2Y��v��8�j������<���3K��Đ���7�*3���F�uR8�6�!%�Ŋ�_e�Ֆ(Cp���_Qfe��F�ŗ�_d^�j�(��%�T��Zw~j�@�)�eh�cl�A�R]`�y{���y�_e����&�8DsF�M�p�N;��B���?*T�mµx�������q@��`ʽ1m%f�1�Y��w �Zo*�4;SH��2_�b�Ck�l���LQ�SfpCg�YŊDV�Ɏ/��;i�a�p�B0�P5��M����(�ldp�#T�#��-zv�A�¸6d,��j�c���Fk�*�M�_�"=�E�-huOK�e��0��m���F㖍L���i-=�N��®}���N�N ���K��)�s������Pyl.�s��cm�E�
�y2�Ɗ��>A�֒x�������I?l@c0��f��
j����)�`��_�G���]�t`f�KB���%��e�h/�%V@�@���=V����JǸb2�2بd��&Y̵�!Xڬ���|�f��ł��U4b��Q�h��H4�XegK�C���U���V�JU�T�b#S�g�^���Q������c5��1
��M#�ʒyk-�K�Lg/�)>w���b�q�fD_=w=`�vh�Æ�&;xC� �X��g��0�r�?e���
��VCSG�.����A_Ɠso�H�v�S�s�K
X�<���=%7�p���O�O֜P�p��k�r�:��=3*��gI6'��R���l�~у>���B<���2�-�pw
:��b��e�(�2�!��Q.�Z}���ܠ��oc��C�?Gs?]��0?#�5j�3�5��r��n���C։��@�H	׏(h�����[4�r���l����q��m6���{Q���G4��Ҝ��PQJ��/�����8tn�M�!S��ٟG���g[���0 �4f��Z�I.�rPM���!�k�t��Y�X�h#D4RID�{yr`~B�ك�D#^�6h,z.QK�K�N��n��@#��	!2x��5	_ш�k�4OuP�4�)��]�r�
漹,�i�i��+����R�n�?�(T`������g5���"����>/(3�:�^��H S.eE���	N��sA��w��><˩mLbB<�@͑������*�gCC�}?�J��s�6�Q����m�r�&v�YX/%Ĝ�A�\���I�^l���p�P�B��K:��������8,�P,���cP�h|��U�R݂)��E�L`�i�X/��e��A�<�z��T"�p�����_.�;h����B�И!�	�עV��j��s���_o���x"��<�Fz��F�G��B����ݼ�kG��He%7|�Y�R���m��r�{��R�o�Z�}YN��Ny��3��}K�Q8A�Ε0Q��~��.�5����Mpji��=������-�{�
�5MM��*o�4-�A�+�Er+��6V����C�O$WB�5`��͑��~�H��B/E�u�c�z{�o����$+��%��-bY�}D@��}2k���衛1�f@�0ߪa���d |kU]��}W4:}L�Ŕ����cN1'�W�R���=Ŵ+�'L�j�� !�-3چi���F�BkpU4ϔ������b9���Q2�	DӮP�B9�����d{]�.�0��78B�ɂQz, �d����m�x�n�q� A���u���r��3H�N���rI�r��
i��o5vE�5֛�'{}msUKqǟ�lX�&�GN��]�j"��g�NAj{�->+Q�U%w�0}��HɸQ�Z�l*�D^��ԡ2��/�Y%�!b�����a�٘I-�@����82J�Q�Y���A��M�S���}��]�������m�����cg�Փ�q�<�J�4�	�0{ ��\�a��C�����y�{����J�,'*��A�v.!���o�6�f4cZ�0`������w�OI%2��
��W��S���DT�T|xu�JQHj��Y�$�.��㛚P�Wo#Z��=����˯�h����T]s���38�Ջ
śF�.���6�>Y�jQ�$N�pf��4���#B�M�:���t3��׀�	j8����t����L]^/A��^9<�l��V�!��ׁD�ܨ���T��(MV�H(T%�+.�]�1;
?f�v�v�4r�"Ϊ�ɑ���DC�9�2�;��,�ixV�s=���Ձ௉9�����Y�f�U^̓A�"�8PM}\�Z7�kWE�B?�E8��.9iݕĪkU*~L�6�v���΅�~�x��:#�Rļc,A�߭Fg~����3���A�AD˹�y���3�iS�.x�-EP�g��EZ�~�Lʉ�]��6��0�Ȁ�K"�;���TB�j�hQ��z� ��G6w�ɍ�F��� � /�!���D�݈^T5U�|nR�/�z2 6��_��J>|�>�5���y&�h�A+)�F�?y5Ł�dO?��ҳ�5��{3)�H}�tI%s�����Doa;.��Okd�f��Pizj�6Q\k�M��Q-%�� ���g�철,�k&��(Gy��+*P!�'�Y��?
LM3܊ۡ���(_�c��ʼ,�%mc�NY����1z��C���c�;���߳�?(;�� ��y_-��FD{�b~<@T#j���� gk���V4f��;Xii!_f���vn�WS=^'�M�p��&cʍT�R����S��kMnE"9R���qf�|�C�,��[�e� Y�;x�r�n�G� ��6(�p��d� ݻy�Iu�@�0��s-vf�3�?����R����5n G#�ݮ�!�i9.�g%V���d &�&5����!^ܱ��&�b<��ɴ���͌a���Q崘Z�)7^i�h���|��I�-�ʞ������F�[�P�%R�^R�&�.ˬ��h�uˀe~u�96��r-�������mQэ��Ţ옱��n2`��P
`��ƀ��t�<e02�Ҍ���j�*;���gi��>/o ��Qql{7\dZ�)�����4�$��>����,���������!g��7��'��`i��Uh^����h�yB�v�{p^]���6�us?2�fG�N�a�c���S�c~�����A����-vSU����f���:�����]���Ѫ� uI���߭7=�RδG�/;k�3��SL0v���gA­�_‪��{*|��n��^�j�O��ds�qfYttx�6� \�KY�K����/3��$m��_�ؑc���eg؅��ebk0{:Hp4�uy��̱at�=K�c'�O�D�v� �[�i�ɘ�B�c.Î���3�u;�X����M%QGO�C�ߴ�
�6�1��3t�dU��W��ͽ�,K� �U/]q�� �~���Z`>�K�(X�5��)l׳0_���!"(ߵ^�$�8g.�0�����2�p���+o��*x_��i��_*��d�dr i��-	�w1 3��?��w
X���� a�gLǚ�5�\'�a%H��)z�)���0�{c��i2�{�<h�(>���F�_)��C���7��WhR���� �b���Q�W�d�9}us���pwzO���[���3��0�ۖ���GKL������;N�1�h�˼}8�M�e�E���-�	�� W�/�փ�؂x�����|�/�O�	J���k�Q����OQ]zr�ӈ���v.m�����8�����	0� �Ϛ=�1^2�!$0�k������_���:BF�'xҊ��g��|�Y����U��u�oG���E b��Vi��3�nݔgൔ��x�b���{Uh�pZ�hE��y��@%���
�A_{e��l���#�@9�ҕ��LY�NDE�G�yf��\D��x.t��K#�3˄ z,g!+YĈ�12��p^��B*A0���R�BU�9Gg�O�B9:���/�q���1A�}Է�H/��Qϸ�����8����H���MTJ���zE�n�m���0�����t��l�0�>Y�Ȍh:�,�b�Q�V��u����Z�VaY6DQ�3[��g>��� H���(�(�Z�b�mL��a��.,�uJ��Ӵj�F�� XX<��8��vk��'�s^���{W4�,s�T+�Js�_�(�W���V�מ��z� qc(ka�{IN@�/��G�q��[~�)k�[}�fH��}PL�v[�!"���n���<;�����H+G�q����cذl�z&<[�Y�p�0�E�d���0cDJ��{�i�uqyh�L�����oy�I��G��"���M)�����s2*�q�L���Z�M�xg�S���?��$�܀[s�}�h�V�َ0�����(�FN~���v��ۆ�D��Ջ5���%�F�{n����JI��Rq�\�������0�xR��S�@;fc�1��0Tl7$�41���ya�f���� ��C�n�Q�Ԉa�xq+���R����(�8��q�5���r�����Q��ډ��Z=�]oUXݸ�Ʀ���43��`��C�)�̇�ݾ�I���7Oĉ1��H�ϘK���r|$�}���@���mP=�<����Q�0�3���#ě���)��p���s̈́���C�z!�LL_ܞ�)s�/�o� �u�Y�%FǀG�OA�����h�p�H���T>�6��-�a��*S�3���<Ԋ��]���Ǜ ji��sw����~�!E��� [{˵���Hۥ,��<"'�Ͽy^��Ӭ^���l=�_���i��<�8{�w��	�s��/��TL�w�b��eg�ʶ�����*��M�AK3wV��G�X�5��,0����6�u�+.�[�?�Oۙ
��{"nԽ�~��W��t��P�� �f� �ga`�v�7�2���9�xk�?!��a�q��1Qq�g3,��k���dA��[���I�Vu�85�J�+t�
�u��YTǙ�Sr��s	T��&Em0�i{.��3T�$U���G�V�qx1�d���D�aԙp���$�s�/ЇΌҕ��$p��Y��}�q朡i\K�v>�8��UR���_p�S��6�gqT1}�Y5����z�\2	��$���Ƅ,����ɲ���3���{��e,l���T��-�d�+hVy���2X=w���H��*��KK����br���̷h�AѺC���o��]�)7���7K�TV�"�Y
�hH��3������˱���j�.W��qL�|{����_�5��Xإ�2��)�hn���aم��'�L�5u��h�j9�Ԥ�@�k������A�Ƀ9f�	�ʊ��Qٻ~�(���[:͢7�����AW���Pitu�m�_j1}�}ф��ʠ"����x��,��B���u]|�����IO�)`��fu�΂ɴ7��(�i^��;8K�#@n��7��ͬ'H<�lJ�����W���r������35*��qw�~*3O�3���&����x'�$����:��T|<�ld�KO�=�vf�)lh�,��EUꤊ�z��N,k��U��&f@�p��(5����9e���5��$����+�.pWsrFI�X�	WW,7�:Nb�������G���a�m��%�^0x��#5r�[b=��&�5u���=��x\��u�8���V
�ƴ=Q� �-"!	��;�t�	B!��k��c����/q%�O��dYɡopJ�l��v�h꒦=Qg���xS��������lA�@����Co����H���%�$}���4�(�����\q�NB���`�af1��A���.�٣s��=<���3�@k���0�~F�2JI=H�g��k���ߋ��y���c���B�]�{�3�2�AfI�S���^r��B_(9�����Xw����*8|Ƥt��K�j���Γ�r��#�읫�h4i�}���'�h�������,���9o9�]s����pe	�-�@%�9`���Ϝb&�0G��'�E2��U�0Wm)G�Pa:'OŻLsPy�7u^�`�C�$�[O��q3:���ĬX:,)⠒�\~n��syprC�T���;g��{��=Wc�]��b>̛V�:�H��oG
��(���'�^_ 6F�Z��<B�m��E�Bq�&�|���3��I)�z���z�9x{���k.��K���Fj�~�8�p����;�kDS7YpCd1���lkL�c3�)kц����M0з��Bc=-U���hb�p|�_M��zo<'m|E"��qz\������r���h}C��R�/��:~z=��([Õ6rK��lQ�ʐ�k��ϱT�c�$XA�e��~�S��Z�`���
b�R�9=#��3HƔ.nO[0��p�31Ol�
>�,�B��D�z� �l�r�r��C�[ޠ�N5����̅2��M�ر%�l�)��g�oD�v���=ڮ��z$��_�E^Bg��+{��L^�U<A�ǂ�K�_�'@h{�{ ��Ia�Ý�'���`�c8�X�h���-˂��uH��������蜄��AR������f�aRac�ivjk��ɏ�{J��2E.�n�sȘ0ʄ����R���=��=���{g�mS�-d#�3����u�]+[���<�+hw��6���,������P�Ҹ\ο";1x$�u~��Ϭ}�������^\L���;���D�Y�E����ϲ�PfFG�Xm�Ы�8q׀/c�����B� ��.,�#+Vm��|�O��0���c3�օ��'��s��� �+�<�+�n��wV�}<��:/2��usy������!5�C�u䓱�M�$4�c�O�
�<���8�wn ��+*=�pPUa}�UX�&^:���O�sĈ]���^�̄��<1<�de�_فn��r�����bUE�l������#4��C����7�-ST?)�G����4��;A�P#��#QjH��3ֹa�
{dCR�m+X��L�:�����ƾ��kS��Fs2&�q��F/e+�x� ���Y�3E��G��˅��r'!T��m�ִ*����7$��Fߐ����@�f�N����M�3�Q��Ǹ�؛���R���&�-��4��O1��"5�W��oUc�s�Q0�2m�S��Gƚkq�CT-��H��\�P�t�Rx�蕅lp�`�|OP�:|�^cwt�w(\E<[�����n��Qe/\H�УK�Ś˫{<u�U��iC�@x �,��j�`�|��[���s#f+�[ـu�Ȑ�d��U����k���3�G�NG�e��OQ�gIe����?�e|9����{>��w{�Y��4rQm$�fL� ��rwx���[�w+{6�V5)ݜ!F��d��p-Ď�@	�����7�r�h�eC�R�n~�� �'�aB��=��Q�C�b�	����izz�R8��s��ձ�t���[�
JF�B|�+!P�vR�i#��Q1R�ٝ7���Č�)�":
�&��(#�h����+�y-������;ё�A�p� +u���*}1a�|A��!�z_�U`�[��{����W����z��c�9D���#6��r��J�W�����z��5�i���B�j��ϭ���L�I�QW��⠮���_��k��P7��e��7��i�_�_$����&��$��Oҏ�t�A�ٱJ'*��n�։��_�����זR�]¹<=��3���Q�Rئ�&�t���ds�I{�d�[Y��Z��BgR�����5C�����-�rF9���ah��Ջ|1G���D�=�m�6^�=#p���җL/	���P��Zo����a�Yx6f`�d���ج��q5n�=d�/�p�U'h��g��RC�{!0(w�weK����r�W&<�Ix�4�=3mR�����Z���S��\hQ���K'Bi��ڟRL]����$MsO�I�2�F�:x�t��}������ oj>/�]D~(Q�@Y�/�'kKT�HkH�(b��y:�_�pC������ �Rmr)����|b�B��|� <^��W?�w�~W���[X��_�/$��՗<
|�>q�P\$�j���}m��s��T�f��Gfհ"���K��H��4Z�؃���f��jr�{���su���U,����N�
������K�y\����є�Zl�$��k|k�T�� ��Ih�d��ᰮ�<��hB���/T�"�]�Ƀ�Ĳ�]�D�D�&s�\�5��}��qPJ �`�»�%
�`:�\�
�ڻu�dV,���\�E�2Z�2puF0���=�(#v*M,U�t"�����[�Y�a���H�����(���Z�&�X��� W0^:���]��R����@Rƍ�ي�{��;t�8���9���A����Df��n��%Ji��K������|�`K���a�i˦f���v��}|-��A��k�Z��}C&4&j�5cql�д�Ŀ$���<�X�>^����SC93.�����_�Ct�j �����3�)kN%�0��T�U�!���K&����;�ף��5&wL�>w�?���|�B�o`��G	pq�!ω��)�>i�#P�7�Հju�o�)���Hiv�9����2xg��4b~��DCf�7����J�-�,Xfi��mD�es��f�r��Xw�����soWM���4_�M�ϊ�!�`��ih��b�p�$��/Q�ض�c�Ggy�b��8az5�,BĂ3�`� �wC�����&����	�\ `-�<�W㰧�L=�<\�f��I���P/߶��}F�����~u b-Y�څ��q�VA�{ꇺ��6�h�u��-M㴮2����r�V�l޴ ����-�-��>é����d�m�p"F���3������6wRx㧣3q��	���jY�\��`oX�KD�(BGܬ���.�+��a �?�5:�����r���ƹ��N��;�h���}3�?T	�ݧ�E'
f��=�_���95�]��A��M0s"	2U����(HSJ������)�|�s����z(�o`��MS�S�+M)&�H٥c�/�$���HE�F���$��*%u�vp���'˙�~:���;��}_N�Jk{�y	hz�ڕu�0˛;�[
��շQ�P���)�P��a��g�8.�Ǔ����pV�ٍ��5��x|��ƥy]��6�9߃��i�%B�Ph(�&�n5yᓋ��H�mlɘc�gLW!) �� U�3�w-#i;��]T����$~N>�VaƐf�/aC�c��:RC��$�D29S�6]ˀ�^���)��͜[Gr�v��1]�\	����=�$e�ݲ��nR�*�6�J���Ͷ�0������$��^h�μ�ۙ��;�E���ܷwI4��`�RC8Ph� �%�<��z�h��1�y����b�۬Cl�җ)}ZMY�~#U��0i��0������m��c���r��4�Ⱦ
}f����M[�**{����dh�` ���+��T���|�1�gj����`����MgvṦ���H��x��z؟_�nxL�m~h������@���xJ�,�C��@8Ϳy���Yk�!I�*ϥ�Z���ID�u.�5�Qo�;�=�d[/��T3o�GsQ}aN�yl3�gW�x&�˾��W7�T�y~t��/����c�Cɘ�*��w�|$��n"���bo������=1?-�z���úQ9�gC������ł������?�]�?���� !����h�-�)O�T�L����H��9�ُ0.��>�)aD����n����mQ�d�|���^�$}��M��p�G e��O4��o��)��jo$|�ȅfǣr���4i�~���m&Y�B�c��C��5ͷ9W��d�WK���nM�U�ɻF�G)6{8	�	<�o��j�P��Z�4�m�ңG�3V� u	���9�åU�FG�:�G�(�,��Q,�U�z���Kv�u޼��a�=�銹{��6!�ڡ�t�C��ީ�e�g|�Z`�mi!�$WF��M'ǆ����2j�8��r����Rn�hk�WR=�����&���b���/;C�I4�R>��[�龿�_Ȓ|�|�ï
~�Fi<����Q�#��S���rv�����-���c2v���W�O�_a?�wO�u��R�Z]zÈ3y`��UG/�'�TJ�u E'��;\�sx���o�cb W�<�ف8��v�f,B�b�f��4ųت�0�K�S�v�KO��M�S�4w�~����{� �B�q���&��!�KP�N�Y�i�1�9n��J3diO�~��7��g��`~k��.B=�M2s�;��vJfl���Y*��⛆ Q�������� ���6gM�gn�(��rh/4C�8#Qf�-/��S�
�aS�5K�`�,���N^Vy��Bl�y;c��
�M�'/8��6���&���[�q\���}�wP1H!*�y闤��-�3�JK�Ht�[˲@N�\��.��\�[y�C�q��K�YfqEx{��E�*TM�*=�n2�F���	N_���J{�u��~,4w�����������}����{e2J��/���8}��ʶ��4>�������A�!��R:�>��wۻ��2�vͳ�+��{����	�D�-�2+�3��A�׿�~��b��U�~�a`}vx��P�(���w��&�]\��9V�܋t����kJ�7A6 �l��u5r�q��W��xd�@��X+�d�@g�}CV��f)w�c��#B�Ĵ5�h~���K� <�h�2YGYʺn!��kP^)�7����0H��u�����ro��M�:��)s��,�ZHO3��O����'�m	�̻k��a�bփ�=B�a��oE��ҢWRA~�Jݬ��A�6�p��|�//?/�L�	)��{x�D�����*ʰIb3K�Z�pP�K"�N��Oj�Дyi��w{�cm:߷���%
�L�y�8jMp�������/�0�j?�Զ��hK�X��g�&��&���h�5cO���]��9���5N�H�G�r���N�����"/rą����VW,���YW��*�Έ�[,qB���8�A�?v>X>���/5۾�~��ݬ� j������~6��
��T�\�ED�n�(��e�MR�͢�C��m�����{�F
ﱺ�on� ���J-�)�ewJ�}���Ƶ��ѕO�|S��v��V��ؕ�܊�M�J:5����0JfW󒛤�!�Cl�,-\fO=��4��� S��;�H�d*�~q��'��Bx���(����>�m��v�j"U+v!�������j�.�>�H��`÷���@#ٌ&KA�sp�"W�{��=�����3��ߝ�6�M)�"�Z��G(%��!�_3��+ϥ�J�-#��]&��=��A`�:�\/Yl�SG���ͫ�"�� 5����e.4*�^ȶ�S��Cs�L/�+�P�@w���@N�P�P]�P�Md¸��%�>�R]�\��]�қ�F��e�m����PzsT��5PN����E�N�ʥ=諑�˂;q���_��`��k�W%E��:��Q�Xfݩym͊�2i<D�k�y�"�?���ރ���v�^U�YW���C� �:�'�C}�o�!T�-c����A���m���k �1E��E�i(Mf���@ƣ2��*Ἦ����QR$�ͬ{�M�|��Z3K����,�T�-ĥ�2ej�������7x��;L,������7\���5��^�Y�5?�2PI�]�&�?��z��s��u�A��2��t��_t/ 4��Q� �� I!8�Ȭ�Bƶ�J������k�eK��"ZЊ�0}Q���b�lI�]�d0.���0$��E&CU��2��I��[��`v!Z�F�Ǟ����k��::�[]?��-5�KN!�[Q�Lݿ�[��6[��nk����ە+ ��-�g_��-����g4�g������xu��Z��`�¢C�J#�I{��`���.�oY ػ�HR�e����*vm�໷q�N&��l�?�~�hB��Qie������m�l�I�g�����֞���~�X�}�t���d�������-�A�4���%Sq�47� M$�'ʓ����#}v�4�ĕ1H��H_��>^���o+��x*I����8õ&.Jo��|i@1g4ʽ�����Vx����vFB�@ɐ�_�+[8b�n��p�!���ٗc��^GN�8H����~4,�����A@x�<5��1�q�z}�Ҙ�*�B��I�bǕvѐv��X��E�K��d�>��s�s9(�uáK��	b��#c|�)3�m�(���S� ���,4�ؕ��	^|�	L���?άiW�nYi�����Iإ�c���r�E�pPð�^�7KO����r��y�t�ůNJ۪�+z@�������vΆp+T��_��g�"��:��Ϊ��D��4ʏ�a�qFM��o��˰T�'��Q����MH��<R*VQ��r��@8��s8�rC���س3Đ�:l�W��
�Ux��/u�3Ǡl
c�i��	�Z���ÿ��@Z+OI����8`6"��o��M��,��v*�ˍ$.v�G����q���eu3+_oġ+�{s��,�!?��N�C��tӍ�n é�9���1n��}���;���>�,��6w+��߁%\�|�w�EK���Z:`}�ԗ�ϼhR�Qr�Ǟ�G=<�=�(�PG ���ٿF{�T)w�{���1V���eഅi��i��llPw J�<ODA�TH����+)ǁ�	��Ξ۹1�3 �K�c��m��ɧb�-�k)���z?�sC���0��
~�g�C��"�d�!P��QLbL7P��'�ۈ&�d���f�}�f{���j�_q�cF_;T$7�xRiֳJ�1l��\pF{��0�_�$`���6�,������#F\@A�|Q�,Kp2�o͡����;g<�5b�k�l$B�(�J�]���-g�'�/��J��1�m��e���wO������`l�Nc�*�x*%j
cUJ�o'>�*3�p�����?��5��½�e �L�z�_4i�f��%4�} �3�)�����
����>c�-��m)T������[v���)�p���&#O�iQ-�77�oaJ�?%'�3��$P�t�ؾ����]v�Uބ"�+
�]�K��;6�L�r�I3����eB��
Ǭ6���R6UӀ���H�C��ǭ�@����X��NJ3�ِ�a:OVd�Uʷ�÷��l�j!F�#�r�h��LCf��a����b9(2_n�E���S˞�X�lˬ1=��{65-s�m�\��W>���0$%���$�Z̊� �z������+Y���t Nz�N�M�S-�/<���d��#m+�ԏ����	B{�'k�~DݿG�Wt��O�����6�C<�ZN�N�L�����y�羬Z��C�����3��F۞�B�{:Wm�9���n��w
aI�z4��m�F/H����r�����Z�<�^��~]�q4vtް�#�����zj��-Ș�y&����D����AQI��K���*aҹp�ӆI��=M��<M�"�859o!G�z�&�f-E���|	�P�i���]C���Bɿ4Q� e�S++�qP�e�_;�VK)r�љ��esKQ�:�A�AA�0���[�C��e�&�z]Ⱥl\����=�MG��J�������J���F���9%�IL���Creq����_nA-+<��ֲ��3�b@Yz�����Iܮ72c��F֒`���ʟ���w�uqT�޴ñ=��<��C�5X���(�y��z�c^�Bx��s�����ל�HwG �k�6���>����S�Rrҭ�*�� �G'�h�a�Uiw�	��,ٞ :ӹ�Ђ���GH�+�g���	}�T��9T��E���%�'�'W��z16F��Jg��(�n]q3�U��K��:K@��M+��ꌭg�=
�7�C��{��	��I�ح�F���@X���Z�R*��������8�Cw*��'G՜&T0�:t�c���a���fK:@���[�4��w����o���g>j¢���YzT���QX9����ΆԆR��-�l8��Q�[{'�no8�t��^sK���M]�oG����!XBI���r�V����A�~���X��S[�J�.ώm���E)x�T[\,��HFM�� �B|�0ڿ�o*t$��r�ƕ�λ�Y��ԂM>��w�G\iY��A���t6ʡ���pu���t��a|�g��6� q�IP���a�/K�9d����FoJ	n�ŭ�k��)�x.@j}��z���Mg���B��5T�K�]�	��A��i� :h�
>�]l�o�r����$N�%B���ӡx���kU���WZ�B�'�"L7hF=�o�],����+�;٨TD��)�.N�ԅ�A��^x����\<�8�] I;�B����ԨG��Q�M�p�Pv�LIP�ķ������n�r	��e�F�B�L���݉T�`k<��Ul��J�,t50�Y�qJ��o��:}���I!f"V#��G��f�Zm����j;���������$]԰�������^\�c�E;+�����>3�O�j6�N��T�:x��a����:N��hb�Jk��;�!���ge��p�A�L��B�GZac�'p�N���~B}��ٔ�IX�C���Pv]��xA�Y�|��U�#BX��F�g�J�h�����}>���^�m�M�H)O�v��qz��<=���/�R�s�)�٨��N��G�f�!�\"�(qQ}��Ǯ� d|"Й�Nn�t��h9B��g���&x�*i0M�
ܰ���+CѸyc`�4?��ܤ��у/�&q����髶�#�ܫ���|�-�(A�}
3�zz�b)XS���8N�ٌ�x��,0Y���ǅ7��Ntj�Z�m��I���sA�T->�Ɔ�>a������"q���@��R�
=#%d���)����e���̏�;#XR#�\]p��Y�f�(w��F��;�M�}[h=��E�)<N�ǷQH�v��b4���B���B�[�ml�޶=�-�Q��uڜ��z���0�a1��i4r*�~�9 �Zj��5��.�ߒFq]~�K����叉W��qwl��3|�i����{����S�Y���_�,��K������`��.T��[�h���+����uȹh�iO�x��ŋ�\�G�(�uѸ�� ��M�4�E�'ϖn�&P�BV�q׷?.;�((�אK����U�b���_�i%cW`��d�9SUQvC�q�Ԙ�t2� ^�;fN�@0O �xW:�Q��*e����f�(J�ɻ��J��ð_YU�A>�X��]��Yn����Izm'��T0}(���h�1S^�*yI̿�'Qj����5!i�Y ��� ��w������)<�b����7��Fo��*k���=S4'��Ɨ���?#�L\��CTض��[Xl�l+Ai�Y���l�s��Vx�ㅥH�U �><��6��W�͙~�z����s�7�L!�%�;�&��v.I�K���ݏ��T����t.��zר���;�����5��󑓉6��>e���w<��5`i�u9!�8DJ�m�,z�U|�4fu��"ä��	nK_��|�Q������3$qj���gme�f{��$i�AN��e��������3��z�u�MC˹e�4�%t���3�@����q��~{��[�D)��T8{�;sRe��&�������:�NV9��f�Mځ�n���XL��(�1o�Ǧ�E�I��E-$�X�wYUۺ��'ʹ����8��Y��y����2�e��d�kߘ����~26	��+%�o4З���!"C�4S��3&���FS��e�	�ܶ~7��Rd����=����~�؊��Г`$䀇:g�.�*�R��)��R �B�'9���,�<� uT�%��c��7S�R�Fc}JP�A#G��a%�0� ����јM?��P3�/�ot�i����ž,��'��uj_�Ϫc+y!��;W���P��H��eZe�vѱ#�bF
��tl�����X��o�����L����B��7Hdt������$z�s�^�V�[Ⱦ29Pn�i^LD6pk��?�~�����K Y�fL1"�H�e�����W�{��`@�h�N�E���k�O�b�w�����-�(����x"�ͪ��4d��㺤�+��sq>����s:C�gbg��t���e�N�����%���w�@<'8m�e�k���M̰?U�μ�Z@����q�3�$yH�9�Ο���}��i��;pq��DH��������qEU�5� �ea���>w]�MޚS	}>Fm9�c�����z��5F�6)���ȿԷ.)�ϰ�����_=�� ��>���5�a�qW.B!ة�.���~�h���Z/\�rB@.ʀ J��Lu������A�v�%�����P�]K< @�5s��O^�h�F99��-֟f����J����&z��D�����t�{f8�P���Ӂ�(�=���n��vj?��N����:����� �(��_��ط¼�[S��?�����)�z
-e�zW��C����"��(ڝ��j�d=)�xH�����{�7��������L۹��Spb(|����3�S��Ĵ���l��p�
N�����u8kb��Fd�&.��NnV&�;�=o�X6�p��)��ԙ���pU�a�U��u۱ë���2.;�7ov����2�\�d\�t��a�����ś(�f��%\%s)���Ȥ�
7ϣ�"ޠǕo��C�b �KT���o@CT���n:�C5fE��r��a)�[�(`hz���jo�Y��Q��#x_'PQh��>�>��FR��@3��@^ �P�p'����R��Z��ߐ%��1���ίL�g���5����b��e��������� ��T.��!)2	N�Y?u�V�*ץ�>�?X",9�a?�(��H��g3csJ0�/�<��	�����6�N���"-���
b"
C[�4��{9��ʘ�}�#�Db�G��z�S~*���*��`��[1�w^¸ɳ�"*d��$jMx��W���8��â��'!9]<ޟx���ҽ��C�@�/�O2���7��@`�n�c~(*b�dC �#o�ջ�յ�����f�ߧ-��cKy���*���}������6Z����hyfIv��o%���L���/�3�Sj�G��3�J��%��on}{���r�;��C�r��G�gI
��Z�1��`b�{�[@��3���#9����Hmw�.l����T�%�~���1)sy����}�^�/���m&���d�m�W�l��p	:bc��&���Ɏ��>ԕ@_l���y?-���HQ0�{2YY�
��는,�^9�:X��zw�K�C� �<�����1����	~�p1�9yA~_`N��:�[�?�9����wYlC�4�:l�B�@����V'Sʠ�&h�[�i.�<_sOA��2X�my�=��Q|-2-:S}�ީ�O8pɃr��;�v���O�^P~���y��)3��]� S�q&9�g\y`����7���H+��, A��/���L'9���lM��!���ͽ7ρ:�&�lH�B���I�F��6��0�E,�2j7�ؚ�~�/��L0-F�d1�K6��e�w�	��В��S��4���<��<ޓ�t7�f��˃裐{�.�^p�un0��b���������Hyn��~��V�"��?XŌ{2��:���9׾mՍ&���1��'��6}�{�!�9/���g��Mdo̙r0*���|������}����贪�ޅ�NX�V�1��`Ԓ�m�8�\J$�7��9�����S���9���nmm!�F�9���脞�ݰ�&���w�y_	��R>%�<Rg�9� }P*I�R�"��P"�pq� �QW��+߸<�66�(��2_S���D�=�� ��AfG���������x�+�9$��U�Q�������W�W\��T1�����%��C�5:�E���gpq�XpTZՆ�C�E��/�ܓ=d�`� ��7]!*{,�m�ӕٓ \a(
�c�"Ws��r_�i~�z�_�� фS���R���8%z� t�y�uS dkm
� \���\̠%�#&Ō͉|&��R�*�OO�,mT��B8�[0,oH=���r?��O0�㱌|�SS��k3�s ��B�>50�D������[l�.�"���Cľ�1Wk[a3��v�J��c�l�-W�G��n��Aw���2�l�r�!����*=w�@�9�E+����4��~F���)l�8��{��b�v���e�.kGX;�����#�8��I- K�̩4wrݔ��m�}���q���D�ؔo~���o�c��m�A��~��
r�NLu�/�M�T״��]��ԦRI��좒Ջ��|�YRkM@��R��5�
�'�~�H����K��uir4�p4>�fW�4ԅ�Ȅ���ら)�6SYN�gGQ�� �b~�����\����&�9����k�
�m����@^���?@�]�%����;p%'
�/�M^cӐTw���`"����(]�7�\�a�֤@����k��-�R}y߹t���q�y}�񡓠����.���N�\���_��}~��z70�J�K�OS�������G��q�^l�#X����v����U��xs�zC�?82Ԣ\,���@v���+�QI���8�b�:��?Y@���� � ��Yh���W�ڜ0#i�y��?�@����xY��Xd�'�mW���w<�*���w�|S�{�b)���7z�3���P�J��Uv��DP�w�؏��G'��_&&����1�����"p�Dg5���<��	��f��ON��v���bPA��hW��O~� ��(�a<d�Pwg��e�zW���@�����jDxX^�����~�/��V�Բ���7������R�c�p�����ATy