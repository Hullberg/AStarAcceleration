��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����yD���*m&Gn�h���U?�l7Us}�q��kn����{��:���4D��:�%V�OVy^ƾ��Ž�+�eƲ���;;�R;3���j9�/��B�)c��@�FU���$	4_S�RIR���c�Ͳ�\�
}�Xpuڪ��V�O�G�~�5�ŵGP:��. &T�
e~����9�'���`èH������d��^��#.�4�b���gTtۡ�iW����Ft���ݥ�:k`�����֕�&^�U����cޙ��ւ�C��C�-S����8��܏��ω��+|I��D<�X��H����_i��Ձ_�T�+Pd`�8�j���AdP��U�=���@c���ƀ�M,
�S[;���E ��-�`>�4)	q�ݑ3��`��uA�
Fx�F���l�̢0��(�ŤldF@Kj�sN����p��:�����	�&#����d��ug�z�/N�S	�ˀ�B]��i�q'l)��4W�@���@1�}�M�@���$����r�'ЏF,%��ͻ��vx�����aO������e*߸��\f5+t�Y���hV0�q�Q���R�k>�T��AF5�Cajs���;�@��0,�FHI6�2W�T�zѝ|��HA���E{2��gh��ˬq|B?~�9D�c� e&@=..A1��U媍���2
�E8%������D>�Rd@�K-*��J�=�(
ïx��s��A'��n�/2Co�X{/ o��y�v,8d����}�B�A�Q��f����(��|������ؗ�=�"���_	���7�����1�1
�_��؉���0N����hR6`(�i�)��2l���%�L��X�D�	qv]��B��5���J6C�ЄL3i >Gp��1E[��E�m@-�xQ+\��S�HU�g�1��ziz��4��T�"�9<°��F�'畟�?��<E�_�19Uz~�BH���K�\H�@�#�~�(x@�� *��(���{�����\h��y�E���\�����Q�����Vm�$u%m2�F�1Ŗ�t�|	��6	�����a�~���W��K�6'S�𥚓T���&?U�3���/*�E+� �~Ķ����\)J�����8���#������F���Y `��@9�
�G�)��
����QT���f�X��!Z-�@W�ي�Bܟ��DQ'\�>�k���;�f�ǿ���6�dZ"Ly4"T?P�%A�4�&s���D��Wƈ�IW���.�LS�Y]5����l._��6hG�B��2�]j8�R�
�'�ҠbY��*�ܐ1dQF�
U�"`i�!\�N|jx=�9Ϡ���}C/���4�Q�k)�-SQ���^>��Z�1IO�:��u ��ߦ!���gO��W��i�v�~��$�L��!^��.�Y9s���J\� l��}M��s��η�X�����$c
�i��6x!ZIe	�q��7��GR��<���-b���d�����O��˚~�<�7p1"�g���&L�kO����G��(���tiM�����20��'<:���|�g�B��S�B�i��u���� U@�i]�I�qU�͊2(.�ͪ�,��9��g�v�3���Wo���T��@�c7�����Ǥ��ϊ�dK]�"���f�b�����A�� L60���V�k�@���"�B>֨@&R��l�k68�l݊3��R���G�uZ�4'���Uʓ�`-�7�3��D]�o�K�O8m���;X�q>��|6���ɘ���٩ﺜ�8ՀT0b?�V�7?��$,}�,b����o�F�xKYC�����Ueb)9����C��8N�9s������;���?�ָ�a3Ihh�앩��h.�#Ӑ���0lk���K���j(p�(�q%�3�X�{�r��a�7�p����.Y���^�_��+�Q|d6:`���rO�_��#1����X#��Aok�p�/���-'��ZY�ů��f���W�Lc��+����-E�j��
�L�u�{��8��j��R`Fow
�Y8"x:O1c]+�6���@��� G@ɮ�z*�ٮ�p�Hk��(=��q���yo>S��"Ɯbe�E��c�
��/�5��yr��e2����J�΋�_�#��^�q���ߦ�C_�m��s������z}ѫ鐿;��W;�lF��*��OZ�EJb@�Qlh/�8�I�oԲ�,G*@8FK:�E��/�)R�x��q������.tW�6���?.�vңK}1�����q�}��nkHy6���onх�dx�ӗI�-�]c��@Q��K �������k�碟FAi,t��M���DOe%o������u��2���dtJhb ��?p`3��W�9@K���uh_��-��������:5�`H.��#�k�Hsdԟ�o^�
�a;6d�d,{<��1��;�$���Loj0��7F���ʕЗ�#g� n��-�yp9�n�k<�l��j�׈ߧ�WC\
�Wox��WZQ�Q���8&�ҵ1��h.X4��@,Ϧ���3}�jA�����h�Q<ؔ5!����r���;]�|h�~y���#ʿq�¯9�׸��X�Svb�D�s�LDO?eEY@x�%.��i���I�ǒRS,��qt���d-��&�W���_�!��&��zIA)>vӢ_^Gjz�y�wm�@A�0�-��9'��*����w'X�,����d����"��Z�3�ØЃo�E߬A�v���F�~����b��YCj���+b�����G���/'�gx��9̦Q1�PQU������q�]i����M��8vf>Ff<[zw�1���N�e���Be��s��x��:��t��c�~#<�������x0��dH�Ҕ\��.�5��3@��}���'�+���L��!'�6��C�0��+��S�$Q�j�Y�ړ��3I2��sCq��~��<�90�%�P
j�h���Ci^<���;��blV�/%:3��}������_��"�i�{����M���ލ\�͔�����c�po"L���)dMj�	A{���f@2@3�w���_w(~�,ɧ���}�1��ی��� �f
d�E�N��.�^�@m��F~`����ұ&��P��>$�8&Ӓ�_� =H��(ϧ_�*W�P�'<�+.L���y/��� ���Aw�6�#�k�B`#��	_�LKG�x��D���87ٻɐ�q�/�=4��t�i��,���s�a���Q�(R.����t���8n���L(oEg��>n�ˉ��:7BM�<�j�������<����yO�_:&$��+�nUy63��t�ly���Λ�ڕ6,ZX�����+�*,�8m��{�[3�3x`d�������+����V����(t���z'&-��?�����e�׆�#,�E
��b-�!�Zl��(/�˃	>r5�&��?>���X�ʶ�e�a�R~Ɲ�|ԏ_�g�Ͻx�J��ڹ�o{���yT��ao�t��@'-e����w�-n&h)��G���?&U�k{/ y�c��	��i{a.�W��`��\�I��ϛ����˸�H�md����0�]}�f��m�D�˔o���*i.(�K,HR��Z���qf��9��/.�lp�[��$���?C�j,��It(B����� e�~�K�[�x�K�pѳ����g��1ŽF=�f�τ1K$��� ���>��7�휧��Iv����5�@�-ż����Bv{X���8a2с&"��Yv,W�?ed��Eٻx��b�.J��ڡ�'Crs!Ǖwl���B4J;$@���bL��*b�70ϼ��RD�ɪ��Ɯ�����RQ?��$� |x�d�.O�z,�5�����>�Z���8&?�k%�\U�;�M���:c_z�"�M{=���!�NCY?���q�e#�eV��q�MT�W-�[��Z6�:�8�+�����4t,�^��s�(u��BE󰾋>|����h:�������܎�e���UN�l���rU����h9�V�+O�V����6ꋾB�D�$\��V3�J9K����H�
��*�0:��f�D�h���Y�n�9�3���g|��̣�+�����G�C8�� ��V� �ip���(���7gM+�w �a�٤��A U�W])��Nȍ$���w�� jW�r�%�~�G�i"����¹�:
��ugG�652_]�1��n"��<�X"����t�q&?O���5�߁�/�TL���S1o�����TbHw�C$����`ve��LG��FM���_{�B���Ȣ[@˓�Q��b:�Q��2�$�2v�dm�ʀ��z�����-v�w+p4��vc3X��gH�+�$}x_/�W�������7ε�sJ���u�nt��G��a�U����r`������F�D�02��9���qM&�6�|��do��eL���!�</$�{|��i7����,Qy�5FvJ�BYѱ�U�n��(�#�	�NQ_��}n��U���E���ϱ��.u��Α[i]�_�,����X��^�ڍ�ŭ�|7�,u����E��b[ȡuzf��G�����������Z]�4�a��k� <�<[�XeZ�!�I���~Ix��$�7Z�w?���6}��U����'��)�Ÿߒ0���|/>8�1:�c#	F���(I�/<��8
Wv��1m߱eC��ېhqK7�5c� ��q[�����,�b�K��ܘ.ܚ����9�(�,��I[A���ڼ�ӳx���^�i�Mf��y���+�ij�5�B����X
�H͐��u�K��ܓt��Z�H ��HJ ���:��,�I�k�����=?*(���^*�3}��I�+�e+`%c�[�O����(jB]4�N������j���z��(w۱�}l�f�����v���tS�ÞT��#���[���>����6�/烁�(�k餚ˆ$-ˀ�q�K�e���ח�".A5�w��f��� ���^a������z�E�ρm�X�ϧ\ru<3��o�|�a��y:��k�&Տ��;������-?+�U�9��dxrL�f�7r�0&��z�eJ��}��Q���9C���Eg��V���mS5\c���eeҫ	���7���"8��Y�h��B֝l��h��*�6N)�����Z���}�� �Ir�št��J"ܹ̋����ov䃟2��Lz[�ik}D���y`�5'�!ٚR2���[�/^�6nlPk��@/P�PE��<	�3u���A�Q��]���7(���۶�����E���YK�`=�>��g,C�i2 �6�,���4>ų�@��$�I,G���&�5Ϙ��:`�G�h� ����=�U�&ކ��( >�(�:����PKT�B��%|��~~�
���~�ci�_p4w7�N�Ԑ�]S:��$p3:�!b���������
���P�~�ߖj^�㺧�Zq"}Q�:�݁?���7l�l���f�8I�m�	���W	���R[�G&x�KK�<F���2� 	5�q�����K�k�?�!R{�f���8-Y^wc�pU:8�Yà�C����zc�}tf��y�"Թ9� z0�{zs�o�r���	,@a�GL�zv��|�p�W��w/��OԢ�ۑ!kb��o.��?%��;k��H��y��a��|����������TI?ǧT��rޗ5<���~U-9-24*up���hO���N�����2�bBVAHa�x`���6`������:�Ŵ%�WFz�]h���h���e��$���FBb�U\��@���7Yq뚷+9����8g�.���$ëa��Y�������_��ID/��Q�����۳x�ũ}�i6kiTЁ�[��E�B��f��DY��
�eņ��?{X�ҷ�V"jN���{����.�D
<Tm**�Ym���_�+8�~p�V�wި��.����CJ碱i8�#�(�S��h.�h8@�
l���r(%��\��Q�$�r����b߱\�h����6w�����FՀѺ4�	��#�~�T7��b��ڋ�