��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!��ߌ�6�u��S�`T
��E�E� -�5x8�ym�7�4�����Ƹ˲[�B�?�O�aT2>v����BL�j��>��D�7�i�9y/�_��N^Xl!����u�l�_S*�
+O��\���~,�Pq���N���zlO�<�/��5���i�f� M$E�wנd�
B�M ygiz�NX���LRg�LGWqd�[��J�8�/rK�vM����J Ŝ�bO�X��r=N&0<=��&cA�q>�d�(����~���tO�_������ȇ}���f�{��,Xh�V*G �r�ܦ�u�V�g�������D�*�d�B�"S��y]M�j�������P���D�E{IƳ�5�k1�&�;��ƨl�A���6�0�
�V������ެ�x�jt�@T\2�/.T��R�헉�q.����-��g8����(�yև�Qn�!��g�L/#�k��@2����dzXP?�p�i5�v��66����9%����vW��&嶑��Л2���;{�>���_����+E9i����
�TK��0�z���2i{�H~^E.�[�Q����q��-�2'v�p>S6��Y��g8�'�\�����Ϸ��Գ�M�]�PO��W]|>R����Ж�������#����������UO[��]��	8��E+�V��9��P�14" 2�ٷ��B��J����H ��@�Z�<��ftCL�Dvvw���,����Q��W$��l�̞����+�)��ݒ�
�R	��n��5<�����&/���t����w���b��Ǥ�-����n?u�6l��H���3I��_� ʃ�V )L��*3�5ַ()L
�����S!�_&u*.����BY��=�AKq�flX�բ���_�L�V$m�6�0'8:��t��1�ڡPS襞Z����N�/����%d���:ҏ��X�a4u����7�^���IS�j��a�A���Tߗ�	��������&g{H���t��*�c0����*?�ܜ[�'��?�t3�k�R ���[���R�)&��dhl�V�G�l"���!N�8Mf�Gx��٢r0SMK�����%�yڂp��y��� G
���j�ZH%����\�{+x��+�E
o�����s��\9�c�xx2�&�����韚�>*�؍��`��/���
f�gon��%���T�}GS�W] �i�)���b���^����Ly�\�i�<�&3p�=�G?��S;�|ڰ�TN ݠ\l;�,&�,~��o�v��z�`��*��W˃�5`nI�d�/.]�[�q�]�g��5f�!�8�nb=��(X2��	*<BG�nuig�+k)t��Sa�Y�JO�W1' p�>�s&��=7fօ����8��֓���{�W׼���V'Ȼ��� mz�P[9]���a����}�-
o�m�?����i">I��C�=>��64�)]z�o	 '��Jnuv�5�e�F�����2>�c~�A��;�e�v@q߁��m��ls��a�c�i�iJh�x�#�)�' H��'3ܿE�؞�@zd�97��r��-�=����X7X��B�y���-����n�����@��T	T֙T)����򔧌h�Ik��˂^�H$A�p�ˏF�����G�R�s����	<����Ҏ�>-Fr]�;(�!ç����7w��O�#({F�E��?�K��O���:sVT���
3ț���`V5L�����N�	���G	 f#�Ηvٹ�T�z
fS��@���f��UN����j��|��Ѧ��Q�Ww�?\���)����F��E>~�-��g�EX,͊��&F�ǣ�RE���r��kGآG�׶b��M�����HW�`����CnAz܀���!�_�B�X4j�J��t�>���U��oj�4���1���%��lto6N��l�g�9����M�u�d$�69q����$?�t�n*w���f4B��G3YI�[�t�������qU��S�׎r;a�S��NwƩ:�/	=@��?֜M(�4@���o�S��#o���4��
7:�)"V��ղ�1�汙�g�Me���W�X��0&}�֭���^S�!�� AsR��d�ь�C��'⓻{�&�6 vL�;yA��;A�"��MtO���7���C�Ռ�/�?i�)�5c�IC)d?�g��p�8ϮC藺Y��,)J����e�}��^3��R��9���,ݰ��|(�v��w]W����N�Oy�欱8��ߞ��̷OEs�د{t�j��\���~%��:K6p��А����qv����L��6��A��S*ժ��)����W���\�}3d��ۀx���3�+�D�u�g���6ȿ�d��E�։=:��X/��[u(jk�i9`��Jw�Aw߁}���ݔKٌϣ�k"��x7���O�����|�i � 3
�a�[�	��l���imZߘ;޸�� *��% ����`O�:�� �C�`�V�ϖ���H���TvP�On � ��H��Q֜�;&���yLvن��x]L���F��"7�kqq�@�:�5� �5�e�:����t-U�Cg����~�΅��#K�����7b��uk�L���^�C#N�J9�^]����A�}�Ӈ��aP���0��*��Vډ�F"�AJ��9��6���Nk o*<��yqN�;VDF֩�[��x�1��D�{�=&Sa����W�����:*��l��ucq�T�� O����'��s��[�`\�԰��-E�h{�K��q[+c&Q����`��E0����"�i��;���%
�&�0h�Ԏcu�uI.�	��a�Rхܗ�5�,7��MϚ�{'�
;�>��a�1m>��T�]�W�p��s���|�~�A�Uz�>�ڪ 60A�!���J���0�?l��7���-�ڊ:P�X���?/	GT�U�pXu��'O~���B4DG�uZI@<^�R���='������!��	��`�l�+$��=���k�W���F�"�蚮�������Ҕ��t'@*��o�΂�%��^|�4k��2��7U��B��t!�)<_zߤ�)��o��_{?N�����6���>�W�| U�wIv@N@#U�����{ �o.1���f4���u��\BslJ'
((O�u�����kSkJ'�:j���ֺ����Fג\�uՍŞr\�7@�Z���Iz�WE�0J����g�;,�T�U�zp��W"����0~ ���$u�;�� �J����Ϸ	�w�P�afe�SQx4;�Ĥ$�%�t�;]��8��i����8q�GT !��.� �d#�Me�i,~/_+5j�@� Sw ��@3G[$��yeJ��5]�<��5D����mx'�����4s"4u���$��)�_�0�u*�)�܈((�����7:j���|?���{&��`�Ny��c���˳g��5���U�m��ՇO#u��u��.�Ό�`[E-A��Q�&��y��S�]�vA��7Tm�hT���G��Y�A}ֽ�SS�jY}p"#�ȬJGH���0�.��bk@b�����P���Թ��WD��ed)��deFrB���t ��7��K�fNƚ�3kw�`["`4��u�3�}����������T&}��P�ֹ�����#���׃z��˚�����$��S��1�J�O:��%� �>ہ^/����O��
�3?`~�V������<�r&[K��}ز]���]t%&o�#\v!�ڍ���Jb�bw�������iI��D�P�E|�sZ��v� j�kt�����@4��8~8c���������8sc��C��ڧܐF���ʹ�^��p��u��0��^g�i�ƶ�F3����'Oc����o��T]��#���[.�"=4j^�P.P`���,oUH�~�Ќ�Ι;3Q[F䙂�Tg�+�Xp�G����z�M�Kq�DG��Y�e�����iN,��	��|�!�I�\]�W�1�F?���<
t�s�t4/��*�u�0�<����n�������OU ���U�d�5�����G�f��G��ٍ��Kp��;�KF�Ir���Q�iZ�8h	�hW5�����UIT�3��#�_lU?�*���9kA���B4_2�
�S�}�=I����w�y.�㝞9���td�Nb���W�,�\�!�2�#MC��3o����(�IsF��ᣲLފ��WL�,��@��'�s�IW���� �K�WX���DG����i���o0��(s���]�7lm�|+%��1������<ŉިB��.gF���#��ɛr��'�^��rK�4˫w�G��7��H��fb���rE����U\𯂩�fW�S��ԃ��'_�OՊ�P�β{�o�Oh�H���������hbBZp�zG9�
m۱I`}�Uė��ʢ��a0���֞w	�d+Z�:�Q�����4�2@�R��Jz�s��_WI�k��Z�7�v��N�O�¸ �א-�s���>�S�xy�����%��m��J&� ���-�A�B�NZ],CW���Iz%C�Y�[9!mܬ$��4�� (a9iiz��1�kg�p%��5E��p���d(}yGfE�mD~�]������?��R�΁���Ӎ��b�R�+W0;���"��� G��D�Y����%���Ϟ'�N�6�'�q��Pqx՘ËԸ1�P�A�j�K���qt��D�(o�#6f3YF��С�{R����g5Қ�Z.B����<"�k��*��폋�y����x�~$f%aӉ�����"�r�z2�n]��=��[A���U,Ʒ�A�	�znE�`��N���3ܽ�u��˙�&W姡��dM�����`�w�\,��Y�Oz���Ri8Io��`�T�$9���z�Mv����z�9�Xfϫ����sS��Voa��ʓ$�A�e�!:jN�ꩦ�K��2�3!��������qF0Qb�A�C�
�¢��m���d�g�	u�n�tg�f
����+d�`��RP��m��ݼ�� �$<�k�\rjӏ�Lz�t�w�1���a���A4MAP	����9�m�>Ctʇpi���c�w��\ �}����n�=��ί��I=�%�+<�H@q�N����{�����A}�YG1]���~-�t�rv�`"��O��{���	�"�q���>q��Z�:kdpk!������2�E&6nW/�ՋD�n���5��0����6s%���%�М���$q��'�H9 ˂��"��I@�tQb���d���lT��� yK�ι�Mm�b��LV*���|��H�"e�x�Ɯ����VVXN���/��Ȅ��G�k�$�e�#i1��'�B���뒀�����v�2�0b��爒�	����t�c��=e'a���T	��w�N��nd��i晝���3��9��H��n�"P�������?��1�bu�=��H��]{���g,�nb�S3�+���f�1 `�����|�+�Ɣ��U�&ѝtsn��l���NF/�+��8!�I����e ڹ�v��̋��ŵjz��YK#�"ӕuNS��1a�W��/d7�����4�� ��O[ޡ#�ib~OVt�yE��7�A:�X�R��� OI��x�r��皤����T�b,�V=
����GIB��q���>c8�M�xo��cǲ<g�F���S��c��tV�К���R����ĕ%��ITč�㫀��ur�\9F��	A����2aM��r�o��ZѬ�������oqs���a����K�xV���H���Ik��t`wϾއ'|�8z.��W�!�gK9�|9r�tHY���S�͇2ɧ����`ؖDO�[{i:�"p �/���X�n+��c�_�xϹ@�d5�
�����uXǨa��)�CE�I%`	γ)p��
�>Sf9ԄVD�T�2����f�of!$��m̻��x��B����X�g����4\,|ؘ(�Pl���e��Q=�p�I�*k�s���XE���\�����X�G
B���I����B�t^��|�G�`�*_
��1��T흐�6&c�0祁Z<�\��<\`�H>���M������9��g\���ˬ%C�J�N(����!0�R��#�R�+�-����;医�;�F�1ЦX��ಈ�w�^K
��h��O�0�cPe��~7�EA6[�PÖ*�>S��ĉ�ࡁ�DU����p�PFkb��%�7��I�A�d�6��*M�$'���t��c>!�b�X��Aj���?�b>����Xn�g����C;_G��Q랆�pToA�K�!��ש"��n�,�K�G+�����68>㦣�@����f���!��!��8�Mq`���:�K�b�X�Zzn��p�����,�Zx>�V���}7#L�Ev������&�l�6`ĵ�	�L���E&_72"ΦJ��~|�/4�Z-F]�
m����d(������2?J�H��8=6�2�3�������'V"r���#�Q�@���r�RX���ߝx�F�����@��t�h��hY��G&�k�W���xۭ{�Z3�wP�}D�J�)�iז���oy#��&���̾�N�	�݉�F�g0 R�*�!J���m?{�l�� ��h��Q���xh��,Yl�¡����a�EŖ6�z�!��vE�?�Q�J��5PX���T0�\39�o"J�-��#xu�e������mcJ�����">�3�c�����\%WRJ'�M�I/�Mr������w����el�N���5�)�?��o��&%dgp��s�P��>��NH(*`y�w��x�h����CO$���M��
���|k|����R�7j�p��4܃ټ���1%�s���%��M�+
VM2W�����U����v[N��atP����������+��x𙈈�������vv�v�b��E4��ۏ>��h�	��q�R)�FZ�F6��U���<J�P��HG�H�u��?����.���"�|!�+��z��'�E݃,��Jk�j�I¢��Ѹ34�ʥ@��t��؎��?�]�q'Z���;�>!�Fb�l-F%�O���v!�[�0�Q�����͕C��g���K�-#V���-#�g�G?�p�����h�ս̲2�諸������aY����7�(�;�2������ʕI�O���@�z������[j�::6%��=Q
��J�'��5s�M��~���eJ'*+ם�����>��Y���hdWo	?Ud������'�A�ۦs�n�MiM;_�n ��a_�N��e��;wۼ0 ',~�]����:�=x����0�����G�ٖ��y���1�	�����̆���*��^,U�"g����,YY䌽:\�7�l�i��rMBߚS��D�����
�=��r��m�����[�����0�$m��;Zl��m;+�m�i�q���$Y���Џֵ.zOI�u��I-ǄYU�vO�e;�Y��ˮ:�.���c&f!9t��u#q�Z8�"y�!C#�� e����}<tg	6�v�W��Л�Y�)7A��QdǺ��dV�I��$h��0�d��J[o�{!�w��c��m�r�� �Fֳ�d9h�MP5GƢv|�� �R�d�=�4�}m Qy1qT��K慴]{�î����%c7�ӿn�5�b���G^��G��k(�T�T�����~3��$�R@��a�����VS��u �>d������c|�r�R��$C$�!L� ����:���a2�Y:&�ad�y��Q�~��b��J9-bf��3���P�ތ�S����y������I���Άl�����.[g{dC>����^Q4�o�'o�>H�h�qq�9�����+M���`������--û�b��lY����ѧ�AT��دB�3�A<e�m�Ss ��`de�5a_)%�>�s�ќʓ�T�Lvb$v%�Im2���,�X�R�p�u��Y�/-Vh�l�ަ:\�G��4C��������l��p�G4.��>l~�"��̕�6�d�SR�R�V�ш��f��Y"��Hs##D� Lq�uv���o+��&Џ"��|]D�4);�J�W�з$�ɐU��r�ܖ�7��_ng�^,��qc20��Ռ���dёĆh�����~3a����[`����h��P��5�*G�Cx���E�b:V{��>�S�����j�P%
������%ʹr��x )� 2)P�s�Hm�-����x�]��:n�^��=C!�}O�# A��V�1q߾<���׼n+��~�\1� ٿSnD�68������3��� �W^3,��;�s��^Y�%	U����h/S��#ҏ��H�u1�8���=?2j�`���'����W��<C
��GR� �w ��?��#N�n�%3�PM�݄\Q��;eGP��y�K��?0T�P�A�-�+�m�i����� ?���Y-~i�e
������ţ��^ .�")�x)+FtH��۰A����}�S�ʿ�Z�.	"L��M����r�+�ꓲ}Q	ʒ�Lg8����.b��{��A-�8dqp�l�� �Mx��/��E�_�%�������ִ�T�r-�⦲�)ja�����@�M��ԛ9n M�$��Cg6:|O�2ŴG�l�8��񰗺��������j���4݈�"�a��MO ��R������R�I7���Ί!�֖�򆥆Ug����(��x��E�Ur��su���ǒ��lU|�^�;����_�e�&��kqSi��͍���'�Ua���WZxKy�N��.D�g`�����ʲ�db���C�r+0��2T���p�5Ŗ�G����:���C�h��� Q��������+��M�3�fy[�Ξ�H�<|3^%�[��f$\���I�4��Nֲ�M���R��SZz1Ƿ�rx%��H+��l�:q���a)t����|��S[&�m���s�����R-�PR����.�;���vX��l���B��aH�l�-�߄+D�bF�n���͓��1�W��]��\��2i�Z��b6j�G*Z����������G�#�
4E6@�a�9�FE9*��_�����U�j�69��ڗ%��Z�)9n�tQ$��j�ܢ�o�Ϟ�W4���{�qKo�+lB�Tτ��D��W�NE9��������w^�t�ЁKeV"Ẏ}��=�$�����&s!�a����P�WvW��B��P�"!�#��DK�c�|����|D��I��=�7�1!n+ͭ��;�%��o�H�\�eD��&F�j���W�Jt���U�o��.��N�:
yn�/��`,A7���H86tWg���uC�q#\��r�g:<�S]�ﾝ��`�.qulӳv�g�̈��(��ڌ���?y��5l���;mh�=1�t}��KI'��$�V:ǴNV:�� �U~ڔ/����,Ef~�&	+�\�'?.LV�+e���������<���2�/���R���L�×RS4�Z�4���y���˗V�� m���f�0���r*���Y�%��������(O�jA��^�v�Z@'T)�Q�%��d�,ؑRj��/�&�e^��y(�6����v���\�rf�H�-=yX�G�/Wf�n�z"�[�ޚ��&Qx�e����˄�D�!���t]�b�iv��f�+>[C�`���Ӧ>��e�|VTm�7.gbl�����`�Ҙ����Ur�	Ĥ��e2=\LMU�DF��*  .�3B�r�^���R[s�6�)�E����s���~9ȱ�0ydE!Qٞ���LFT�B������wS�kVD6��;.��,�7U�D�.��ʩ)����O���Ao*b��DAD�ܠ��ý}������`G�7]�t(n��������)��x�
�N��Ѯ*�^<�MB7%O&kq׸ϭ�8"#�Xt����Ei���}�h4N:)>�/,t_@� �XLΊ%at�˛�*�n��ϔ�k�6�/����}�Y&s�Ճ61�E �pS������]�B�9��'�4�|��?*�؞�v�_�H�b�'�3�P�0�WM]m�T��� x7_�$�n�2�)Q/iu(6�5�C�Z�?c`¨�f�|�b���w�b�o�[��W��4��ܴ'�o�8g����&&[2Bq:�O����D�T������TEe��"�^����]&�K�q|'>�Dȸ�"}JIX"�5w��Bm!r����k:���RI�<l�J:�s�Ib	#����KOJ��5��%l�{gxO�`k���j����x\��G���">���L�-n�}�?+,
X=��Yz~H8+uN;]Ӊ�5$��wM8�A ���c���B;oAhq�N��Q+ǒ,{V`��b|������p�8?Ol/k	�d�|���@>(;��z���L�D����<nϸ��2�#���*=�t�����K������R�T��Zw!��8} 
<y]a�D+�bT_�i~�ņ���t��,�6����ɦ��̧�����kt{إ<�Ѵ�q�,��W���_b"7ɜo��l�7�im��4`S�Y�p���?�_�<��]5,��%,V���$�[��cQ-�~���-��d� ����{�A������M�� NM�/�mGh�řE��i��z`��O�/K�s����pe2�E|R�W�O��뮮��Om�@*��UZ5�B��W���2R����X'E(u�)�ɄI�����K�p��s�=kUaZ콖��֋�3�;��czTQ�|"�V�n���-Ӂr_�ܡ��t�F�f q7�8�f����nM��%YM�;/EP����Q	���t{vx#9�V�h3����I�|8b�J�)�?yS`ښ��8��F�F�^6yˀ��67�S���PJ,d��I�Y�Шo�z:�H�4[��¸9 �6�9�Kڳ��ƈ�I{�s&`��'[�cN,�C�~�Z`�Ŗ-������x/�CU>�^�h�q���èrǖ�5�*�j]����	��P����[_��Ly���s�3��O�E���[�&������DI���`�w�e�1�cd�P��	��������
��=y�W�HT��m��=`mF�[�8�X`k�����qV���8�)U�7\[��L�9ɹ�y*A��r��`�~���D�����BJ�� co�pۀ����D%�a^s�	��M����.װ��|!I`	Ѷ^���`tTd��(��M��Q������%Y�+�Y����Y�n�8�X~	��A�b��D�ȍ�[I '��V�8L'*��ļ�;K&�F�]���	b[b|����*^�"�(^��0��7�' �m9T�>Ҕټ�AgBiH
��߷����j�G��,�I�C ��&�t��d�D�p�0LM���������?\t�g��WL����D0^��v�F�\Ui�N���8�Y�c�x�d��vඕy�(_P�n)�nt�b%+Z�VGPr�t}>�3]ӱ ���5l�tG:�me�����)�N���a(!�t��[�g��jx,���p#=>�g��w�>�'�$�8FDy��i����y��"��9�;�d&Ŵ�o�'2h��T}쨩��mł}��hH`f��g"��HP�9<�oL�:�p������󇷛���W�:���}p���M#�Vi0�R����?��A-"�UjSL�#O���m�i��c6��A"���{�Wf�1���3;�	wp��מZ����I�N�"�N$��wkW���C,�������ͭ��D�s��xT�:Q���k�oVw6 ���h{���W����{�q V]H�!v��oE����D�VGT|������g;R4"�q�y߂O��}��r��e��Fu��&�6�䐴i�<5F���S=O��H�~�P�0��g��U�� 5��ef�y]y8�a#�����Ө���]�e����|�w7(jCd�h3d�%���3�ǚس�х��7�+�gg�$@ȩg �&���<d�YQ��G�u�Q�>�	��}�`�'9��:��{Lf5�@�����]���ˎh״�~�/�
�i�ƥU�$L1n�\�#�(�0���	PfTżJC`F���_���V���L�������������'@��.&��:,���M�.�d�m��.ߙ_�S�mh�;4x��YR�
�<���)������d�Rz�U�f�P�נ���&i)�N7�Q�.��x�jZq45��f�)�+����=����?���iGj3Z^� _��V�I�ΐ��T���IZu�&�>�����޶Y_�h'�����?�mi��bR0n�5��6_�����1�Qi塪&�\5��k,�E�ˮ�y�d6b���o'�y������:༳��j�ѰISu�dC\q��d�z3_���&��gօ���G/@��%�v0�7̾�o�7��r�ޝ����M<8!�c�a��灠6MvZ� Z�g���'�-������p�n��q�����|�nqa��H Ȇ,��OT�����'���Ծގͮ} {��w��Y+���y9�y�"����5j� ̤��J����)j��O޴�ܳ��M�K���f]�:~9���6(�T�/���ţ�bz!4l�KPWϘɔ,l�lgf-�(G���}{ҡ����%�=P�<�g=pwm=<ȟ�[ޟxG&�J��IA�߽��4@�y���μ�`��6���ز�n��ɩ�+�-H��;����2�J��]c�oR�HAu���>~��d���#��+�URa9e&�ꦤ�D���k�!
>��Ƶ�
Pc�V`4�	�ʭ�^+�V�����_�hE9*��hO>t�i����A�/��bd�*�u�*���� �m7�ج
�!F$Ft>+tN�+�#F�}|"(w�'�-+�0e`Z����a_M.p�p,��Ō�Mh����� �ɏ��:�{��m�����M!!���㗭Ql���C(�4�r)v=F:b���5�܊��Ăbc�fGb���x0V�o޵-�SI�l�4�sP�Y4u�$5gBS¹x��mMJ�h�C�[��W򥽀y��dHꁔ1��6����9�7�KMj�;��Op�
��m2x嗸S�6�O�y���2��IBu���ф�)L�pe�Kv/�~��36%w�y��f��w7�� ]���iC�J�}x	C��p���o~��zq��U�k�9�ez�a9c�d����g+q�/Gb��a��2i�Rf��[��9��z�g��P��6���D�D��*VWM����ŗ䑼ub�	�ʈ�e
�3͜R�H7K�Z�X?%-T��N��l?�eGJv 4v:�8�+�9NI�;hA��fm�;�#�?z�~�s����~�1�߉-\��+�u��v��v�e�J��{aR�Nc���Ȱ͈D0ea�R�\��X�Y��M-��M�ɸ������Ϟ�2�{k��]��j���@���<�,CBԧ�����|d*�z��+�f�����.X�4�>�+'�GL�\O�x5�'&�^�SA��
�!=�<Z"��,QܮH���s��}�'v�md2 ����Z�{/�Mz隒��4ew_�茺�1}`�gh���.�|����
�����+`$n,�d�%T<e2O���C�"����L?AJ���>X�`��A��:�����D�{�I��^o�1�7ҥ�!�}��T_��Z�B�B��>-��؈�~�R�h�2є���M�g�T��볆��K+#f���á1hlOS_{e��~+�RZ�� ��n&�LR�n�uc����Dg{eIg��%<���)�>��3� ��yQ4�ޡ~m�e��>�3�Ic�A2+���r��?�B��w�v�&Y��M�Oh�k���[|ڴ��N��`�8�����*�R��E"X��y|
�lW�P�����dށZ���xCaZ�׽��=5�s�����H�Sh؛��F����4�	�B����ܸ�QzW[#�-Q�E�]3M?za��+��fV.�#�������/����<�܄�ݗ14�`9e���bQ
�s�-V�WY&�]Gn��E�5uҵ�M�LW�~)3�7�Ѡ+o���j@�z��3 ���f�X� ��<����=��\A&\���C2�-�����8�f��vm���pa b����kƨ��Yd4�3�G��e���6\/�����h���s��z����#��O��� ���7�/���Uc�< ���1��8:{ω8�~r-X�2���i(w�rd�	k;;ꐲ_a�0����s�{� h��]˃`qF��zEM���U�ţ�~����τg8�d3��Gu�j���m�#�����ڀ�Tkmj�+�J~Q-�?�|�1�����1rK��ͧ(��zF�~(b�`�uhb�`�����f���	J��^�6F��:/U�YڭOI�.�����w��E( ·[?�d����A*�σ�5�	�zl8�� e?/}mR4k�N	ʚ-XM/Y9Ł37�?�v0��|.�Eǲ�tmܾ�E��-�H�>�����儠�,B��e*�5d����L�
6π��[�:۟8~�-Qv��+�����w���GS�"{���꧖��E�����2k`�}		��Tn�1���ۣ�))�o�k��t��E�N�����������~}2���y\�:?�欭S߲����_I)�hk��@�����~�ڝ �l���+b̂à1nwX݉�q`QGuA��n��Է��� �Ҏ<j��{�}9�;��M�Z~5�3����p�g��8q�!!W4Ζ�G�������{�>*&�i�,����r�f�abdr����{:�<��N��U	f�`	Ee��w/Vt&�X]�8�� �L6B�L��m�P��t�?cr<�-�	��a\���J���T�H�Υ����\�z�+�u���a�5��*7j7��a"=���Kޫ�,�4���A�E)���<��}RVE�%	���ʂǆr�q{����2�1}�����s�ܞ#V��H���R�)uV.�VF�Ơ���%��|��w������$ıN�#0�*�x[w�fO��x/�R)Kf�7��N��u�2-.��l[J���De(4r��B��b��w�q$l�8�p8(5ϓiX9�H���s`�|���d:�P)���a o\��y�Yh7�:.=�&7Y�m��.�v�q��p�	7�8'a�|���:�S��UK�_�4U�R���si,�:����.�H�e�5��M����L3!�k}/����~�1թ����N�GǓ��Z���պU�%ٓ~􏃱!�Hh�1���&�,���\���-m/x+���#ŝ�wG#�C]���?��1��{�Zfq�ΟB�II^#RwzI���@��U��Ŧ�-�#���0![�S�����C�G���ق8��)N	dv2U�厢ռ�D�Km7Pq����r0�2����	n�aP#��*���bN��Vw&::��L��5ŸhC�#:����Z��$�����4��F)�^�����H����F1�/<��]`B���Á���KJL��Lb�i(ٵ��׸c�������n�Ȯ���5©ֆ�����l����O�H�Y:v`��ng���ߊ��=�HQ��^��4�t}A��1������'���>�H�Չq�ߜ�]��_l�a�
�����k����	X��2�]����l�%�d�8�M��U�(�ѿ�Q�&��;W�m\��T+CR��?5v��86�֣ cq}�ۃ�R��oA�-��JD*k_����D<��2$�.������bn�C�ѯ^X�6����#�IAƁ(%�B��]Ķ:����g�Kɬ	Ʀi?�h-�-M;�^�`��ב����*�1��v�Ź"��+����ک�w�h�4y�=~2�+u��u��Ð�T�8�X!�ل�7,�<;+����22p=p�
/�j��������5s_ր0������{gI-'�=���K:��b� ~�	���yKj+��ߪ�w���g�HyN:ɔE�ό�r�����z��b�*��&֍8�'�v_�U�5�RÙ�������]�U^Q1�& �[�<���c�w-O��<�m��	��!*�n��I���[b��3�R�O����~t]/~R�
%�s�g5m����5���:��3_"��Cm泭��`��"nI1
2����\��j>Duy�nB<����4
�*x�"za���z���C���ׇEey�9_&��"-\%P�����7�f��b�YP�M�7��=�Qx�Ƹ��R�b����el辐�1�MjX)r˂����
�;d`�Ȁ��J�]o7�mZ�Ǘ�ļ�2v��6j�7b�3
h��bc��)�_n7�U�����mI�a��$�&tѸ�d����4����M��[��]D�B�7��EE[U�W�&p'�|��4������W���b���8d���D��<k? pX��A�r�;;�� �p�k�Þ�GV�Y���bg�
8� T�e�����i܊[��.�p�2�ʴ㫮צ��ė��0Пމ_�.o����n����2�s�H�l�_�[�g��6?Ix�?~��,�řB��:��6gm�\�B����U�o9��8��s�2r˭�P|��I\2F(Z��x��?���G�:��"���7WF����F�f8A�b]�|��8,y�6�
(���=/�2�dT���M@��������
?I�@�W�W$��]v�q�j:�I�}��ΞzM-���M�t<��rX�B�W��@e[�Y��H�V�j�bpҠ� �գ�t2��@j,<�*yE����N	n�.���E�|j�m�D��H4�{��BDZ�����B�Mu4T�����P�li@�mi�P�z	P����&����|�
���<JR\�(xF�|�X�-<rˡ�;>8(*=��s'��Q>����R]��%a`F�����6ф%�d`��o�Ui�K�I�O�q>�K��]�P{�W��H"���o�m�9��~P�Ƹo�y�X��&i��_�l���|A�W#z�����  �����Mۇv�g��9�DNE�{��S�HJ�)���n�j����b�"=h��x=d/� �EA=x@�>+ڱɅ1Z�Wl���d[Vlҹ�<�e*�(��8�o��R�d��W�ǁ��V�|,\��
�퓃�������Ҡ�Ʈ?�?"x2xm,������������=�f5/4��Ҧ?����2�gJD�I�1Q?�#�A-��]��4ha�C��o��~���2��'��X�w�f;.M@�e،O��3���o�-��;�+�!����3���T���B���2�+�ćL[�{�h5MzU����	W���6�j�1�0�MU�'������Sp%�.�L-p"U߳���O/�7z�3h�B��w8	�PNd/������-�r��ju���ܯ6�Bo�~����U�WPY�-Cw�ˎ?07�Q�y��/��9d�w�ߩZ5��H�v�.�v���A�@̙~T�N��'m2k�ɉD/C�*\�#~^��������	�sߨ�Vu+�1��8v⹑�F��Ӻ�r���њF$<����W�t�j:�}���3:�&�8����G+U,f'��ߩ��@_%���Er�P�R��g��2~�st3RRۯ] �����Q��u��p��c-6��{�ٝ:�9��d+%�&W*5���l q"�}&�CPZ�S����H�O�4���[HkQ�@W�_,>r��-I`)X��J����,˲?�a�Y��bvP\A��U���X]��"�&g@��`Ӫ*�F����>���acc�_�����;�a��b8dM�-���h�z��I�<��F�Q]��>,������ľ��^W,�,��t�U�����A�w2�8:c�9k���t�Eߝ����H���VI�1��XcR�6�$���ۇ�%}9l��Xa�C�-<�&�op�q5��,�F8��xk,���� �v�O$���J}4`�eߣZ qf��O�qv�Is{7D����'��]"�#�����qw�^��RvGMNH�(��O��K��W�W�&�5��k��F�����.�FH#R������ek:�Ӡs���>��ݛӌ�~4�5��'46�>P��L6]A��u��ܚZ�pYH�*i@�X�S3��!%)S�!�g�Ɔ�*��qX���͎0[ӹz��K��f�`�;���h�`.�2�x�I5S�Ӛ��C���q�0�ȬO ?��k�u���53�;C�\��"��J=�vg1|fK�0(�Y�s+� #�L<���[�X}U�V68�JDtq$�n_WN?)q��H���6�1�s2i���U=�C_�	坎-2T�D���õ�8�1��].8������>Fh�v���!^���o<P���ĸ@ub$���'���7��C��PQ�O��绊F0�3�� Y�K㗶FT7\γ.0[S�T�=V��.�߻`(��Q����
q�R�}8=�g���ʺ��/K�5�u���!�Z$'щ�'�4����ME�56$#ʖ��Rx��%�l�@�^'� 1,�l��-�|w��5Ӄ�Ire����IMv��C���xm�ĝ�!ń2����Uj ���&���:ή�=P���{�FVy@���"K���m���T��ٗ����M,��amO+@�^{Yu6>��S��'|�g�8�l���I���ϸ�8ͻ)�D#W�U��w��֮��x�!���DWr��  }f���Z�pp���1�H�+h&�t�f懐��dY���^e���Tr&v~��=�-��s�(����s�R ��F��h�W�Y������ݍ�uE-���7b���� ?V�C)�l���x������bqm�Ӈ�y~f*m�E����/Ʋeq�g�3�d���A���~C$^��$nϺ
�zjd�A�X����,��D��8:5��n?;D`�ڲfZ\ݶ�{g3%���.Gб���Z`�wN�۾G���\3��@���f�}�4�ʂ!�>���[��-V&~���R�R,���޻�6ǋJ�|������8�Î��"��h�)�ۤC��C�ٳJ�����1,�`�k��{�e���8"�W��v�t���Tz���S#�H�!9j�C G���e1T��������z�� ����2��1�gu^���0�(�27�q�2g7���o�J��_30<x�ӹxҧǾ֗��q����e�n-���@�V�[F�@����~5T`ф���t�f$ᣦ�r,�� ����s}�nb����o�Xs��Q�R���=#h�B؜L/������T�H�N�~r��#��q�t�\0vW�2#Q�T3cOc���=�,�w#P:f��rE���W�p�T���z��IBL�������
��������\���
A�5�o��.�P����kG�O�03(²s����,�|LS
�5�О*$�b�l$�n���6m���h-�x�X�'j���4�7ն���;��~�8�ҫ!�1�H�%�������1P_�F 2�rﺑ��M�$��t�;��p1C�S�ity��TQe���r�fى!ᘩ{��` `ǅ��@���UߘÇ��%l=����ͲD�9)��_S!(wN[5j�Q�EsPJ?��j[u\��3���3U��zb	iXM$�	�}`�L��N��"~��U���%����zc���w��5���1��0!V�} 76������aB(���g:����T ]?�F�@H@�坮۷���>�����~+�/.{R��t��צ�Ow �:א�a�I��We��`z�A>�>'c�x�mr6��Jnڜ8Fd9�����[	���\ߔ�˛�Aa>���b˕���z�B���r8���QmZ���/,�ݵ K�ު���ѤkÙ�X�6�Gw��/��)��AB�^W���
ڶu��"�tf\�Rq�i"�g�rT���E��)
F����T�X��÷�oj����������AR�F��d{F����LϺ͕�g;�-o��Aj7]{�"8�"�i��n�����A��-�j3���g�х�� �ݷ(�$|����L6`k��`{�Rw�q;Ǝ�eo��)n<�-�z�7Bgg��9�^/����$\��x>��sY���h�}Ⳗ|/�d0l�Tc*� [y�`<H���N�h�gjLAP�-8EJ7���=Ж�i��r�^�s������?��3�[ ��ff�:SR�P9�޴S�I*�!N��.t�7�r�z�|��8A��7Υ�"
u\p\��=�^#����[S��H �|��#�3��;	X�RԀ�3s� {p"��6�O}��R0�F�w�vp��;?*b���58+�Z�#�a3���AC@}�N���U9wޘ,~��$����]uDQ�,��b7��"�R���f�ae�J�"g��Z��4�S��Ǔ���0PS�\��a5���&{�,�6ǠEl���/�U��k'�J��R��00�|��[ڋi��6Ī�f�eߜdBcޏ�h(ޓb����G�(�լG��;�d�G�@#oz%�Y�y;�UF�Ŝ�BL����~$G�(��k����O	�jz�����[N��O��wJ��a	_�G�G�.>��.��`ˢ �;_��^i�u)�w�,;��崹��y�<�_�S}����2�y�?Mm�o�(m��G�
�nD���H�2��p�Y��Q�3ɍל�n�����^�/q~O��$Ry�`>�J1QI>v:�e�Jest�ͤ�_J���H�~R������H�������42��S�J�'�z�gm�Unh����,�a��{����Pi8h�{_߰X��G��۪]����f�����/<���x��u�
0
9�-"�A�)�_P|����С1`��1$��8���?�[��4#rT����h��l�x�^�9�w[�]�@�ﾎ���|Tױ�z�`�����rE�t�jG�q�9-���*����5���V��(��L�<�� ����e�j��}���3(�`�H{��I�Ŧ�3|�e�s0	��mQ�G��0�!�� 9���f�ˀlW�W8_������Z��sy'T��ǋD���?))):��A|Ӗ�f��H��n$JԱ���--f�(�3N�M-�����F�������o��l(p�,��Ҏ�u��O��o��ٮ�뎭�$v�*�,��(+�����HJ��N�)�P�����CM7?3R��t�_�����UB4�-t.�	_���A�&�ý��q�NMߕ���F��i��qA�BMY&�u��h�j`����|hf�"IA�=�ޕ
�O|��hU�75r~<f�]��f�~z�߻C�՝�غ�Z�Y�6�mg�\�{������8G���2n�^)�v�=�@��v�0��A�ր,��W5�()���N;n��.��rXrJ��	�Il%�'�i���6;�����q��eYh�.s�h�/�t,�ݠ�3���d���X�O�}b�bo����;�3_����Yi��N�)W�-%�?�JI��fAzvd'a�Pn��
z82���%Ҽ.�ܵr�5����s0�?�t�&�衷w�>��yK�̧p��-u�cn�)]t�\C�F��9�i� �7���i�2Y|4g�^�0O��ֈ7 ��;�0���� q�����J�Y��Ȃm���j��$}�÷��v8sOG<I[G��\�ۂΰ�c��2M���W$��3��bĒ��*�o�y.����f�d䦠��
���x�b�ɖ��U�Y����$����=τ-�ĥ%���?ۅ�\�P�&�%]�C�&����S�>ѧh��@m�f bݷ/2z�0�� ����:��)d�@ե/��E �y�,��R���GH��_��^�s\���j�|���2ȊP�s3�
	��D��x!����5H1 HK��@�C�b���S��b��S�����\"�@:���������%��};-��a��u|��I������7�;�-�C��F͖'2 Xܪ+=*����> ��:������:O�uA-�b0xZ
w�D�"��ߚ#���5��n�"�R�O�qEH�*Uvb��(?��(�������2 ܻ		�M>�#:�3v�"MX���Vv��хZ��˳������� ��\݀�P)q�����2�> ��(�a�FyY�vz�R]��Bb��3N���'i��%`�?[A�⚇�ٵB�.�%��z�����UԨ�������@K��w�n̗� ��n�S���$������9�kK�<2(z���q������XdA��������h^��z�Z�7q&�q�߉3��©�#�:a@��yp���A2�q�Z��=�2=m���5�5m��ƪ���U�����I��0>�Q�'�Bi�����4�������+�ff�*���LTb�J�!X��u0D�HH��S�, #!Ys��@P���}���iF9�JTj�-��+TIcQ�/��������iR�dņD���n��p�<%[$�Ŏփ�&-=�loumn�$�g*8�E�D\0�Nȱ|8�g�}�N9@�/{��_������Th4�&b�&+9�|Z9��IZcb�C��&�D��=�u���MbZPY|ǁ���;�yf2�aO;�>nK�}���J��������04�S0�
�k�Ѻ���?~H���D���XEM�Ei�cc���5�Xr�q���&��R��9�(�,�z���=Ϋ"��'�j��:��Ľ��q���L�𛶯���J_��t��vG{��}ʺ�!�1	,�,����W��6mΞ{JJD ����*�	i{���x����(u'�,3��F�,5�_\:&��"��x`@k�0�4R0Deο)��&?i$%#G2ⱍaɟ�����
Xxa����[e��R^g�/f��������5��aQ�J���yk#1��0�f!m������ve��v���XvH�9\���!�__Wp�{�����'�f@ Ƣ��A'V �Z��s����$�n}6��8�g϶�K�Y���hK�ݭ	�|+-��u��9�d�y����f�F /����/��K �x�����I?_��j�~����Y�f�6��饡-�c���Ǧ,��xA��'$ð*��|�uZ%}��=ĮU%�ٺ|����CT\�~ӯ��i!ٞ��M����#��)���͆�Ý��(�����G���@��N`o��W+ ���_���\�����~C��i'C����� Q��b�X�N�wu���Qp�h��R�3�2z��%
�hӸeWOa���l�s�[���3�
A3o����؍�&uB����X??����(>g�%�D�����dŕ���3�CR=���&��;�����w%��N���eFt��0�$���ь�/Ej�@��  ���<�JNS��8KN����>�wRF�ՠGɠ��`23ɰ8���Ǽ�k�&l�.�,aE�dVVA�����G�Tn)�`xwn0��WɌ�`�( �	��/�*�QS{:�ߜ|�����Nv�|�`�P�	�]�Yp�7,մR�>tq|,F.<,A<<��ʳ�M������e�y¬F�<�g&:��v��~�䔰 �"0�F-�BKcn�
��[D�[�9��^o� ��,ޫ����?�D���Y8>�����Nt�N�p��:��t|��^���e9?�*���>L�>��P��'������4����@wՁ�bP�ƩVߪ�`'��W�u��\�w�r�nCQ�`�WgHr�����'h�G��n����v)�A��#�A��x�����8;��2z����9�N8�z�D��r�rof"��#	��U�����r�M�L�'��c(CV=�pޏ^��m�
��a>SO��a�m��Cn7��X}�q��O��?&!O��]�`9D�F���	��η��=�M$3��an�,b�$�2��
Ax�S��v=q���W5��HHù�qܯ}���X�4Q��HR��O���^����44��C2�k��e��21�ž�"�H&���Bs%ʂKk2"@�2� H������3�hF4���k�d���@k��W�����든�s>_T ���d,V�"����"��+M%�1���F��	���mb)�H���_o��C$�X�	���y�����pYk�5s�A#*q��h�U(�y`9B�m��N�m�rv�[�H����P��e�ˌ�6���WQ���(:4�E!þ��.��s�mtc�����;��2����xR�����U�'�!3 iV �E���މ�]�����b���@�m�>�+������k ��x�6�<�s�tejG��g&T���n~z�'�,�e&��+��Q!��cU�XsۄMS}MX$�k&�0�~`?4j�V4��D��	�;�o%�+ʗ��0k�79�Ooc��q��������qY�������z�����.χ�&��0� ���tۿ�>�{�D:cHԟ��?�x�]H��@���$;$���B�
x�+�M���l/˯���M�]z�������AC��R�M��j�%?'Z�ۈ^��<%��]_�QV��E����X��l\Qc	���'6n�PIQ�gȢ2�������~��P���`���X�U�G�\����A��.���*�����	�?���L������>`3�x���L�[�jӀ0L-�J����h�P�&��-HM�lbr�L����n�H{g1oĎ��J��&��DVh�>�ώ�}
<C�S�cSl[�p�v�f��<�{3E���@��;=v�4�8K�z����1�#�{t��=3�>*^�I� �L�T��;�����"v�:�Zg pfL@��[9vmϪ[}�?mrV@*�ND]�`�?'�t0n�I{!�����pI|�8qB�8��1�}H����Hg칅}���[�lITP3�ya#�I���&�]Px��,�2�%�K�w�������%�Jz��V�j���T���źq�-d���x��y����,�� �Vu7�-���!7\ ��^>h�U�[U b>�!j�E�ge�!�f�V���?~%��;��~?֣�R�F��um�Q�T�p��|)���:�q�P,4��p�J6���7��Y���c$C�� A��np�3v���!bޑ�y��;������/!����w�>B?�W�ET<�T��j\gQ>p�\M>X�
2��P)�K���s �:o�]��S"K�X�<��|����~'$����~�j��9��IZv] U��]�N08GLì>چxܧ�;�(�I��GedS`��S#��&���!U�������^�A������L	Z�G�cW!�^~<��5ʯ	�«��4��9\�a��e��pM����G�ўb��~�ۨ�M��/�*�\�Њ�$��\����@�5��Z�!J��ˎ���%|M�v3lF2�toG�[ZOB?�8�i6�a�PnZ\��� ��XD�o1�GY�&�C��H�)��bF�{��L3$Fkj�nk��%Y���n!����Е��ٓ���^�'��+��� !���A�=�k���i��p������Q��*�M���57pu�M��r�����$�ӑ�&�Y�M��4�b���������sh�Z� � �!1)�7���gƖh����?j�,�� ��r�gM�yc���\�VQ�C�	��v\��Pk�C���m��$ny�����}�y��z��'��=J�J\Q1tQeK��;�O~���������10$q����K���ŋ�!0W�������4GS�x?�'(�c.�N!h�D>�,h�h+��<�f6u8�s1=���� �ND��'�_KtN3�¯�[���P�]0�0�n��� ����r��V�~E�;ȿ��R��/�w��Ȟ�̃fVT'ë��u��ĕv�ME͋�T�4C� ��趝��8�ZT�����L]yfiz\��� ���A���V��8�ʿ��5�
0��kѨ�ۓ�M�ѫ,�V�{M��E;���N�L_��b��Ѩ#(�a+_L�^���X^2C���hG�J���g
|LeA=�C���i����?s��=9z=����e��sK�8���&