��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!��ߌ�6�u��S�`T
��E�E� -�5x8�ym�7�4�����Ƹ˲[�B�?�O�aw~��{ᝩ���\�H�2'_�Ь��N%><�Jbl_D{���a��PW+g�:h�`y���1���`�Ik��bB ���Xq�o�����B/�3� O!�7�Tef-F�L$�8��ymVp݂��ʦ!|��P�U��fέ�5#ј��qH���`��o�G���F�?
d�p�@�Z}v�÷Tu�l�o�>9���(fv�'4���".�������9KO�9��KЙ�C�#�//�K��b].1�јv\�	0F�d�xD�a9�O�k��ʲ�=ZH}�M�A���q����>�Fm�-[�-o=~\nZ�����Xv�xWM����폲k�1!��cg��*�b ��>K���Qv�鈡'�*��\�ľn2/��ޤ&xi�N�p�6l�@��ß�I����Z�̿�t6l���b�e�>�������#\T��������h��=wPd��W�aچ"r��]�����K�����o���H�T5�&˻]�럣8��n{�m)�yf��C{O�;� Z,(��/>�ɝ��qO�[�Z�/e.9��2~�w�`6��S��Þ��
�$F�#/�D.g�qai�(�]7�� ����i�{P�fl��<�:@������^8�ˉ*�_�T�5MP9�tX
i���qpb�pE�λ�x�0��|\@����2��b������I[G_"sP�&��gJܹz��h��@�j�{AR86���}N9tQ����Ϸ�	���o���c��B�D�_��G��mB�lQnj�˱����������I��nD�ɺ���G4K�E.�ܧ���fM����+���-�j��u���_tq���Ħp.�������8d��xi���*�&���J�gEV[s�1����EZ�f�S�<�����N�	't���)f%��٘QB5��vU�`=��}-��
�{v �b����4�O,�RMg��G���%Δ�����0@p���5;�F�sB��4��d�İ�;�;_^b}����岩��|���V:�l����?�s�$I'�B�}�h���&ᗜ\�0�'����4��Q�L�����"��w���6*��-�S���w��f����<=�&�T�ZI���g;
�/k�X�'�OH5�i��.{�b�T�!Z_�u7/��0ژ%�w"�H#{!�,���*�W��bu��˯[٥�'�O.�����g��<��}�� �#��L7���Y}�!�رw\K�X�v9{�7����XH�~ 4�W�y���EѶ�<��?�/9�05I�OXv�1.����V_*s�+`d��N�H�ᦌ�X�J�����t��'x�J��7��h�k�NAy�`U!.�h>k�Y�BL66.6�9����)�X�
����QZ���X0����{��#s@�Jg��ŧ�������U�9�����	-�P�5��y F�G!�ȳ,��z)��T�s۩�:9� �5E�}�͵ē�=[��S[��� �%�[�gh�X���H�Y�'� >b�S��v���]'���Xo��r����G���?A��I�V�W��@V�\��&��w�-�̔�P)>B��������?˻�8��- �xZ��#���{F���h,٬{	�jS�Ӷ���~%�t��犺	����⒫j��57hW���%g�����F�)4�j�k�XU��C�;)�k0&c��8&+�h���2�:�2�p[J�Y�M���@ ���:/���iV�a���n_p2�J�)M@J��B|e3����˔L�;����r�� ��a���GsoPP*8צ��l��A�����.�q9:OJ�L ������Q+�aU�_cm��@k?��Q.���{��,vpN�������>�)�j�+�M�Uq�d#��~ل�rԅ��[x��bϱ Nm���m�cT�����54�j�湏��y!��JR�T�Q���R>Z-�F�a�F+�k��u�)Cn��d�J�d�[��j�p�R 2�2�_�"֨���h߫�+�0��`��E�A��)9�? ��~�8�.��̶��{��$.�q��X����s����I%�m�'��G&�H��- �7c6���mE`�L�SO��8܏�0Z
$Y�8�J����BsGF���1�H�򬚽/�y�y~�CO]��N\���(�=
�ʈf��U.Z�|S/���=Z�2PS�X�`b�TP��侲k�چu�%��R� �$m�AQ�2~BV�<{0^n�����uG&Dû|�;��K�l[t��8C~�^��?�Q���}^��PCQ�a���84�r���,�#x���+~ o������_�k�ݔ���m��Q�ٜ������ !���)�Q��<Ry���P0���i=^��dhzo�S����N@��Y��w#.q��7��[�����=G��k��H��~
�.0/��J\�ߨ���MjjWR�EZ��uK�����c6����+�^&�,�)���L<���3u$��<��a�6pX9��X���Vi�h�q�&z�n��OL�R���>*��ʈ�[�r��l��c��p9��?�"u[��qlP����$4�I{�|����?Kwᙟ�e��~�J�x`|u<$Gmt#��qȌ2�R��q�<��Poʤ�8�m#Wj����[5��X���"�l'�0�S��[K͠Y���0@%^���:�H�h��b]�d$+z���Ngp�:��'jw�xX�E�/�~z��e��"^j�a(mF��QBg8]��=����y��zW��F	�({(�#j��X��������Z�1TB��LTw`��μ_Ii2����yCQ�"�MVUꡫ��.T
�v,��=�wD#��T�����j��_#�F$Q@d%)c=j3&D��є���n
t��S�/�J.C��5#��<⮉5ݗW>��3��-
�mb����B�"	>��d��h�[MJq�t$]�AG����E���p�;�/�
�7��!���}Ǆ�Z���o�Z�ߨB���#�&tr�n���#�HV�e���@�$�'y�"g�W@ry��ܠ=V����(K;����%��|����U}�$�ur�'��|Bçx]Z�V^Ż���&�[R�I=��Y�"�d"=S(rn�M ��\�&4{X��m8���]���-�xd�N���W��ug�p\I1�.QHz,���u|q��D�|؋�6��!ݟc�q�]����OVk�_AqȬ�+�$mTV����;)�2�(�|��<��]�o{�r�N����7�������ةh�����:�UY�h������S�4�K�l�k{a��n�R{e)��xfn٫|-t���N/�.q�TSΦ����O���*���zE����
fM���s��o�,��ڭhk�FEs-�t�`�`:E�+,��6'�0\mF��声��큆+spIu�ɇ�+�;4�t�V���+Z�gh�T�]��o��1$c[���(&K@݄%͌N�sJ9b��ÁS��ߺP��6s�mj���<.�P�\(�"WMDp5K��Ǫ��'���H����z
էFyQW@7Z|nD��Q�t�G5����X\+�Q�I�|�C8Ҝ9iW���ɹ��maFvT��85Z���`r�W�5��7���y^�hD4�K�^����S�zB��{o��w�cAM�r�b�*LB�C��	e���F���<ֈ����v�k��Bl̓���&?w��{��#j�� �XDW+N?���x62ң�~��kn�W��S��%����M�ׄ�ϛ����Ho�j�V�L���]����5���;�\f�ޜ�l��$�;yx��}Ӱ:phO����E/8i����[���~�C?$��$Χ�D�58o������'���r#T��7���H/z����� ?�����Toa�@��>[��V�7�A!�ܒ�� ��3�`���%v�� ��m$���aaaQ��8y������� �úk]2��fg4k?�$k�5�_s����H:�m����t^�Ϻ�9���)<�QMc�^06��2��A��{�h,�7�?VH�C��2X�"t��)�hu)��1�"_h�K6><)tv�oq	��=k���|�~��kŜh�-������BS8"�Or����U���TĊ��.C� ԈKZ�*G�-
h��%�'?�	�@ɧ����5U�&�W�* c3
ǗK.��w�h�p_�����J�uc)���d��Kk$p^���a��V�y�Krl`"�yU�%����b�l	Pωw��V7���em~T���е��.!O���ɏH�媤�1g�M�|�D�s���$$Д1�)a$�L�xl��pcp�g��p���B������*�2��N.�$fj'�}��1Z&KŏR����phB�cnȜj@���m����l�e�i��$0��c�Xcʔ2d:���|��	�����[ ?#M�D�z�"�`y��25�p�m�0��(�@Ks�-�)Y+ʀw�@��b��:H�k���G5^�X+LO����m�8@+��b�#i�p��,m�b6>ڢ��J%j�:=:
�Ѱ�x��k_�3U10��w�������uW��=[�^��\k2s�d���~|��5���$�9ug�%�������h����l���*�^��c@2�:�2g]��a��K}%`�f޺��7�bG`�&�������M�n����(Z�T���{��O�A�D�HZ�
�V���4�bК:X���4��e �*w����Z�ӲPhŻȼH�{������xg�u�rm�B�1p{Y�qd�>v	��Y
���1o�3;�.���pL�T��������NR��7�������4���� D�r��)K\�'lS�U��GS��ȝ�4�O��1#���8ס�n�(���+1F�Ai���/�v��#�N��0�c�/�x�Si�(�	���GC��"��sh�Lu1�QP3�Om�kJo42R��(,�9��q\��kc�BV*���dk^�|��B`a/�J-Ċ�,Q�����y�*b����8)z���)��I��N�S��[Z)c�`FVg����?�s�ȗ��l�+:���j��X,t�=Y�C�� QO��Q�,�,�8��fu��k���.�?�d���wa���J0�����~ܺ`��hœ��hm��V���˲�f�C+�	�L����G]��Ml0(��F��WM?42��KOc^���m��r�W-;���a��HW�+��Ek��LM����!�A��D��?��Gh��k���=zx�{f����Me.���\��
ֿ��݃Zs�tN�U(Sw�i��V��9˴�mGA�XM�>�v'��T�S_��J|.�)�ڼL�?���t��N����J*�zc������\�U5'ln���&D��Yst�Log�BV��C�v��\���{<���aK��`���b	�h��t뵲&��h���z�����X١Z?44ٽ2z���l�Ϭ��4�SZu��
s���(���4}�x�v����g?���{tj��e��N�P�Y(%�ȦG�5n�+/j%"4�UR�UE�,���
��0�=*(�rq�<\�����3��c,�5�W�'��Y�#ʼ��>���q���z�ԉ$�|DSJ֠\jZ���,��/� *ъSVL,s"���1ѱ6�K_��:]b�*���*.���r_��s��`�G�{8L���Il���?�^�W�y��7a��f��#�Y릊[̰��&��@������T�Ys����9�!��R���Lu�R=��u��<Q�ql�tp�f�O��9��`�J�he�W2��X�N�'^D�U�Q��|լ�w�L�6M
\cdYސ�{��6�Z�5�����p�r9J�pR��@�w�vbs�@�Z��q������`&�N����=�֥�訠������Q��R��]���C�?��w��͇GcZ*��MRܜ�C)�������p��jG����ƭf�vB�RRn�κ�^*���; r�A{XiUcìS[���m���)At�j�J�$k�f�р.�k�!�{�z���fx��@7-<v&N��������oe�4
�V�L�-f�L��N��jƚ���J�|B�T��Bu�Q�Zz� %��rz��Ё�1���뾎J�]�.�iP�Gإ�m�.���<F�w