��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���q�����W�E�9 Vοօ�̷�S�;(B�����",�U�s����6���i	t̂9։l���kܹ/cFf��@u<�XQ5�"�Ņ,����O��Nj}U��n�" W�u���+F�j&c�l?>"�M/E~�ldPn)b�:�`��WЅ��d��* 	�̰�Z_�f�b�i0��F״NQ�/�3����H�E2l�B�<**�t�ك�{g�9����dH>�7��-�w��7�6M���&@���^�ĔС�m�E�t5���=jj�IeZ��K��*m�@/�L�-T�e��B��۟J����н˷h��}�qA��YQq2���d�4����	����Q��q���W��Bw�^�JWΌ��h3�e4< E�(�(�)�%�C�'W�@"�S��
�Q���/0���O�j���E���N	q��j�ٿ�_�}�o���=d����?($�5�.�e����� kgUDi ��f# �)A��&�gk�b/ڐq�G�Ӗ�2��.C�ۚߟ��f��>'���"�S>k�J�!�I��B֕i؃�?��]��gT�H�]GCa�O��5x�W�wkzYk�;�Ҡ�^��Ϣ�����oĴo92m��ǜ4��q�c{L�F��<v�G��R�����Çj�{�D�E<�~�=�IgP�\eN��H�^@~��xKPWQ~�嵘S/E�qy�J��Ff�3�s Q�9 ��m-�������S΁0{����Lm˺�RCo�gt�xF�I?0���t#�f׬uR��"�GMS�E'2	j�A�4�(n��TWbL�W�/&�.0��GJqOZ;�[��+��s���P�I�Uo�#���b=�8/������H�[�%����b��a�zQ�7n�	�]�2��*��.�����њ$����s����L��1�/Q�V����V�{4ߕL��
�������8wr붐��#�m*��<@Fę�ijqcVC�]�g�ʕ��l��&��r�%rR�Ȓ����{a�~H5ׁ�>���������W��_9ɩz����$#@���G=��)2睽��4\H:a�c�?l�z��qq���:^�Ko�4��n�׏�x͵��p�n S�ς�7"�c�Q�,�RN6����'o,��R��W;�s��3�ዌC���+���h�INѦ+]9�U�/pM}!�� g�����`��b�y�������N!�Q� �}����{-�6)����m��[�`�m���ݓ�C�c��4([R�)�W�`�X�d�ýͳ���<g
> k|���]��m]��M]������������D�}��z`+�1��=:���U{�~IU���S�I�yŔ��&D�j���ā�z�O���^�d0�Ȕ����uA�5�5�bh�r�N7u&���`/������(��#8mw��ثu5�?=�6�Jm��x+���_����Ȑ^���UF.�lQ)���w^U۬��Ν�
$�r�>�=�h��͵J���C_�̷l� u3���q�6�z �7�f�B����T�~܊�D�߀��!�K�\
�S�aXȹ��"�+��m�J\�20	�GK��pL�.�-`p6��U��5A2s^;אڅ�|���('A?.G�W��P�s��W6�D�M��}�1�C�Q[e��&w��0j���'��Va�t1�t_���M���g���F��C�[��&���l��\�x�ٖ��^�y������9����j4,�^�Ջhڻ�'�`�	T��9f�*�)��EQ�TR",y�wW�*S�&V�:��J��2�PtD�+�>|B�p�O���I�_w��J����
V���	��-:`�Y$<���]���Α_霴�j�]��]{����.-��&���:��7b.;�G����Z0��Ǜ��c(On�eV����4�܅Nb����0ށ���,r�K.�z��L��ϭ�H�u��\�7l��<&�#2�sD(k�I�t�XH�='��(���s� ̇y^&�z1R�o���"LFA��^۠ G�P�S��Y���6����r";$��{}��i�MAؓ�N������P����쉃�0�o�c}Z2Ox4��!�h���<e��k30���%�:���j��9�l��f���R��b�qAbw.�
�)���z��$圓(�OG�A�RI1]�G[~�%4���� gu�?9/�g��S]�V_���"����7���S�y�L��#��_%��%e���Uǆ%E���K]�����˅��[RX�<�>/nF�T�	����h��N��P4��1����lJ�AZ� �k �È�Od�shp��e���{����]�~/���ק�-�<W��i�\h��9�vdNK`gn���c�"�dw�k i�BB�fo�H �L˴�K������oB�<2���;�ȄQ����݋&_�_8�5V:`)A8�h�a�ώ�=�bϓ������w�*	<�s�u�m-�����9:��>�j�qW�x~��\.�*X�6�J|	����GF�`��G� ];t�5��Ϙu�$���L��+�#C�ܱ�x��z�g
�YG��N�c�&H�Ŭ[,+f�A�[.)��f`Ip9�Փ/M�
0���A���,^�!�_f<�@q�~��	P��P�F<�`���U�ytB�&'���fW��I��le��D% ��4��!��w��Ĺ4U�7\t�%��;�bWj���u���4Kڿ�v�������ce���8ހz����g+�[�˸��k�&���8�r��tj >1��1.'.�:R���'���yZ�ao�{x0g��5 *vJ�)�<�����Q�l����L����eɶb`��ͤNM�u���=��