��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���qm,e9��Աuű��f�!�R�E�<ȡMHG�R���l�k1q.����QNuRU"+�A�u��4�ZFu����9 ����#C�1N�n\�%�nf��\u�'�<�\6�s�w����xI�H��Y8�/�:��wYɁ�x%>F�?ɜ�1��%��^�|�T%��jq!Sl- B;ԣܗ^E&����:��Y�����^���>��eC1���Þ�sK����N���*IY*�4�׸�?�xh:�x+d���Lp��3i/S^Q�<�����G��6j�����2a\d����e��!�U��K|�C���q�Z�����A�������DV��N��N����i����_J����6=nk�O"���0|�U����]�t��ʆ�\9��1)��y�OB[�`QΓxj)�����/?Sp�`�_\�u��?�ηi�]5b����>X���H��]�o�[h�V��w��gҙ�xy������̹��a�kK��e���:�K��aOnu��k�eFK�O��M�H�H\c�#�X��R0�X���}.�$^S5Anb���c�=u[��g'�|`/��Y�[͎��m^]o�2��f9��p��!!U����UJiƂ9G���?Yw)�bB�}ݟ���:j:���8R~'Y7�p}X�\���/�V*�~����cb�_E:a't��h;��lM��+�%`��1(pZ����3`
CĳYJI������M�B�(!�~J�0�w'��weʢ�Z:.�@�*�pA�L�6��FYЮ��k^"������~���n�Ys��~'��
�ݴ�i�$�[�KX!�`8���)ϗLM�-�{Nڎ��"��6���\���<4v:xx���0�y	fQ�)<�g0��xJ�|<A��!0-�&�*�*�I([of�:�,��70Ąǝ�X^�M�!"@�S(�"˘EӒII;��lXfU�B-�9,��W�|�A"�B�4{}n���l���s�/�tbc�k���3�b]���>��g<8x>$yX�Ҹx��4D��a(�Bꤱ^�fэ�0<�[��Z �b�'�k��S��}�[������m�#�,9������h���O���4�Ѕ����CDe��q�}����+�M�����߅��
�Ie�֔yA���%�cτ٫��ѱ���׈�b�oʙ�My\�%�}��BS�Y��`���/j�G�	K�|'O����Sp�pʃC�u_���Z�����W�]��v:�7߻Hت��P%֡1�?�n��^���c>�501uv���N���-�s Ki�M�;�5�
+��q��"K���ۃ�m�Ǌg%ʔn���G���t�U�������M'�����D��3����e�!���		�])(�E~9� 7���r}�eL��&�VeX���r	�ēv�(��:f�{ݾ��]�a-$��Bl�r��/��d�j����+�oE#ۋ���8C� B+y��
�l	9o�3f���g������`qw��6�S�.{��g�:$��sV�H*=�?O/���RÍ��K:�&{�N�=O�ܺQ�nR�9k%��ȧȰ�u�#Q�sG~;�D��;ȖţT�$�G5'ER<�
;�lؙ��,%�h�Z1�5�S�����6*�~�g~�޾��*+b��u�� ����}��%5�?��� �
��s�	�	���RH��N�qf�%�/��J�`��vH��~$�9�O�9eԻ��~[t��%8�x>yK�b!�ɷm�!����%Z�T���>�v�6�]�a��w���h��ŇV��MEm�x4�xD�-��p�ʷ�y>7
�F��'�8� ��L���VdpCA��!{������� �s�c
n|�����pL�9����>{�"U��͚��8`/��=�	�/S3��;5�����{�^��6S@X��k9x��	�s�z�/#>���xK;>}�� $gH՛����ׄ�U>���L�K!�;�Du�.�Z?��Rh&���
F��Y��k�����;6(�0y�v��h4Ly%��?�o
�j!�`�!��Y�2 E��2B. �I�Q���\i���	�?R���)����k�G�B���0��8��f�����ԆP,��}m<V��,�$ȍ��/����3�{\Ēݬ�cL8�4�o�_�t�����:f�L)l'��9` T��#�<�*�0�/���Gs�sLr,!R1��Q�x�_�¡Z��=W��#�rX�����)�*�^+��6��H�E�`�|���,����U�������1~ �vS�ol���a��{��E��;T1���?�E[<L�#b0��3:ޛӈ��y|��v��K�ꉆ�zW�J7����Vʐjm��2�S��1�/���u[���
!1��ܾ�b��Y�H��^+1�����~:D���͔-��K}�=_�%c��+v|��C���W,b�}�t�K��OZN��Y�ݮ%����y��s����M�{ T����a���L^+B�Uln�2V����N��d5ۓ��p��{*7)�|)Ҙk��Y�R����L��@q�?:��6AIW}��fd���7��X�cs/�Zq�/b���Ӻ3���9
ب���zH@��GZ�5z��.v��ΦF'E�Q�6�����D ��0��ܿ�1�2_��`�^}3��_B���r;x'덺��{D!m	FG�xl�Pu̾n�k�]���k�F�5E�*@��^�I5��ָ:PMO��}���a�w9�CJ��TĲ���R�?�Q������pY�Z�
g	ׇ�4�l����ڢ�K�;'�XgR�SO��[T�(/?B�x�+��O�P@F����n�~L�|��6y�A�?�po8|� �T䅱y��U�Dmx\�'�% t�L�j���gIp�j���Y��S��>	��/���������nQ��\슽���q��3'l� m�&(7�n�JII��[ӵ���y���	᧝��e ��F���dI�*�'�=��k�&\�f��zϊ�&)�!�� �״�� ��0]e����������8�І6P�9���~R�מ757yC�ҠNZ`�������	�gK}�����F�i��78LI>�b5�In'��P�/�CG��idA����j�=���},⼍��o""w�F�Y��aOG�gD���&'���H!W��<b2�~N`�T~�P��{�=�)�\Zͱ�?���)�S�~gKs�^����39�Y|Z��=؉���v�!��g-��%/@�1)M�1������Yw�|��q��b�L:!����6^rQ���9��'~ʿ�] ��� �X�7D�@��г���~��f�@Yn04+^��0R��lE�\Ε�[P�D{[��	w�ӼOa��>Bn�]��n��M��<��缰f�lu"^��P&����zPci�Qo��>�LK6�cx��>�u̡�\�� dh&�l}�E'x�ǰ�o���ȗ��ᠰ��� �|=p�n��߳	���W~f�\gdZUZw+~o1T5$�#�?)�ٿ��GZ�E��J<#[��0�⚇c� =Z���y������	�r�T���m$�z��x��Z��������X������V|�e������9�',�5�0L���9�f�P�>�3����.*L�H5��u��A��?'��sAn)PO��������_vS�1�Ϲ��.�I�v��,3��}�9�`����M�Nb�Eiz�íL0-�,ɞ���܇Č�F�,'3�K7�Sn�D%�JJ=E�/ã�TK�$����Ձ%�_���h��-�𶎽%W�d���[j	P�gU�.�ި^��:�I���,�3 n
��^w㎢"1��I�JQtcJ!FNz�ᢧ3��#���va&K�[��阱�	��("��-s�^�Q�%���]��R
�\��1�}wf[K��^Eֹ�?��(.E�[�	�W%��4R�9q��L͒L[���q�~�Z�i��.�A'�kRW�R�`ܰ`�����6���c���m���Dg#�\\IO~�B$��g�)��	aNVZ�M�E��)�=~Q�cuH�����9 (��;y�~85�Ր�X�1�qU劊�����s\�V�\$�ζp��3L1��4�������Js���#���fq+�=:�\���#ɜq�K��ZƢo-:�I���2?���@�؉(���Ϫ��+���>d��ԾzQ��ڛ�jJ��ZPEZ�����\lIi���c3���fT��8�fO���4[�룰juRw�IR���Z�P�T|�
)���r�{�c��5�A��]��ˁ0H���UZ ����܋Bp����J����3{�f:����o*8�w�!��D..e~Mۼ?VLP�H�%97��@:����t��L1c�?�$s-�E�/�Ԃ�m� 	�c"��$Pе����nF����]�u�o�'�h�]�uG5YZ�+�e'Q�b��X�S�:_#�
�p��ɢJk~�<������?��@A���po	C�3���t������2�YL)!��{��&���"��=������{��'��˟<N(�PLLM�yj:������	��C3���0|�ş��(3�k��a�g�vc���E�ch,c��7ʆQlf�r�PL�,<Uٹ�᥋a��b�������h�]"�a�'�����r�(Y�����!�*���hM�}�%rX�e�Z`�w�M�e�x�|�hĉ�,�ER��t��Z-q�}���W��BϷF#��n���V��6��/�[R,VnK�����C\���:��gv�:]�]G�:HE���l1򛖸ct-{r{b�|0�ͪ��~�Q�N�ǹ+UB��_�r�s%�U��HG��/&��!R��f?!Z��;���z��{����ŵ��dH� 1'��Jn.ۑ�	΂��U�BS���3M���ΗZ'�lj�d��IUV��*�<��*ɹ�����Xk��g%B���5�b�|>�u$Ͽ�6?�I�q2Ǚ��bUƏ�Ӄ �鍋�����'�G����dXݸ�L+�S��$=st��q��"����F�x,���W�VB�)�4Ƅ�q{�L4O�īQ��Tσr"*�wCVC�J�y��y�ؑ5��LD:4���OF��3'�33���CwaK� �*���U�����X��>�X8�|�1Vj�����b��:Yɛ�~��%P� �3�HPT��>%=��Q�rmSe��0�E�CT��##RyĚ���|ݬX���7�1�ȜcȼT��黮�ծz烜E��5�h��9d\A���B�&ޓ��wQrz\?�<�xdkc��h��c��A��mE���wxl9���N@�2P��ƕ�-�a
�B�+)8Q�5�|��*�dch�ʼ�l� �݌7���#p#W�>�A��@��<}�Ə�4Q��D�E��R����]8�!�Ϸ[�Y*�JchB��R[��=zj�}%�sW�c
\"+}E#S���S-�����;�DwF�ŗ����+��/�_ܛ����Q�~Uq�z��[��Kl7�S�~IT��1�	l�'�� _���,A�v�WF��(V�,�)ҭQ�?��h(�F��Ra����Z����T����ؘ��yɥ�D�\�ɜŹ&@���&bX�b�l2��Vμ�W�d�����p3�?sgpz�n��ʵ.__�7�)�������k�զܨݿo,_����j����G����dK���&����"R���,��u���f*��w�B~ ��[����'h�>�LRR1��ʲ��r�|ͬ�9 B������%���a�	���E�p�Q���⴨�(#�RD��s��iK�����7�RJn��8�.�D���4���%w;���y�w��0&Ffj�!ܧs}���\�{�;���FWO���7��d�
3MP��M���<޴�Ȉذ�,RzpÁ�gl�W���Z	���>�!��	7)������~1KDj�o�1#0L�BM���y!VA�]"�����H�6�����a�9Έ�Oܦ��>��h��J�<ˡī�Uq�F�$��S�d~a91I�ڿ!�H;��yg_ȁ�����߇њ���wv�C��=
����LѮ��1e�'BϷئݯ����˃%Qf�;��b��Fp�P҄^0n,�i�q88�{�H̒4(FZ��|#ܲ[�CPr���E��"M��Ő~p�'��P>Mϸ�J�aG;���te���:>L��땲�+(e��n�՝j�z��(�Q�-=Z��ݸd�E�-KȄ3ؕ'�_�=��M�\��s/����r�8 ��v���$�B�~R/"`I���oB��-�X��X����c�}msY����s����(�� 9�ȫXW�^`�o	;��� +6�_��m�;^���v�J�bmz:�j�Z)R�7?A �W�~�%�Kз��є��j����a��9mP놳f�������t3T �eۜ��QZ�ggR�0�ͺ<(��Z����ɴ �§r!���\��!ͩ��@��qu������Y5�:�W�]k�3Ї�w�vɰ���e��=�S�Q�lS�HPk���na��m@���fAZ����h��ژV��O襲/'�3��;L\
@�P���
٬q��F��F��F$�ԋ `5�V�w�Vd���*��y4��r��)1� u����r�y�6ɣ+�Ǜ׭ʷ�^��P�����`��a@bN�������!�%�������o��ߔ� ��;8e�-���҄�}�:�L��d0�"�j�[�R��jz3K�#:Z^�h�j�EL�{�FZ�y�P�~5��v��p��'D��O�L��
�|�!�O<�J*�OA��x��4�ux�`v��j�o?���� �]��f����O�*�z{5��[A�Q�%f���N�s�?�񑦛��<��ҟ�HH?J�\W]�d`D���[MwTQ㶠�P�i����i;�-@]��3��Hv*ҁѫc/�Ka���	���]Z��S۳-��-o�l��8��hNm�b���0@}���۱�ԫGd!����0'�`(/�RG=!��;š�;�Fb䙪��c��pD}m�)�>����ZC��n�C9�U�����̴6���YO�)�eo� �rZ';F�����>b�3ZcB���� �F�z�c����b��t�
�ȁ�*���������}m7sDZZR���R�R�:��f[�?C�d\M�wh�/�
w([�:{�E�ޘ��8�S�Ȋ�6�K��t�h�b����&���MR7�"qZ�o�{��.Bt�NHТNe(DDj�ĵB�U:�E<D�Fgk�u�5��_�j�0�6"�f��}�����gΎk��zwᶫDĨ��p��+�Mil�ؗjJ.�S�69y�F��2_��h2�i�>6QD��^K؁�F&`�vz��P��qqs�{#pW%��*���SϒYju�\b�Y��X�N�A���>R�[��$��\M�v��H�Z�
��e��ܯvӻ�,���:�`�)��{����R=�ƕ��X�W5�$��Q����;S,]C
�Be�r<5�VP���>ߘ8i�w�V`rpY��,-4B�w�hݘ�ip4��� �K��I׏�U��2�q���^5�e�E��8n�O��B��ȕT]]�� �3�\��1[�,�\+�sȠ����x��l}7��Q"����r�f�k���0Dr������}��ry�A,�ԑ�/�	�5� �j%���jŻba ���3BU�}�����Z�}l�v|^׼��'���G�[�B^qI_	�)�4O��t͎ϧ�H_�!�B���}Zr_��e�0�僿 �����-r��%�3��eihj����z�)��-x�]�(�Qʷ:6�{��^kng���:W2��JaM���TU������D�|*|��GA��6��+Q$�
t%��o&��f�q
ճ����J,J4I0�"g֫����L���[R3F�<� �Cr��1����-^Lf,���[�j���jhu��UO�+�I�;�P����Bɤ�>}C��~����q�֏y�Pe�و�z�:7F�̻�P
H���/���vA3�H2�tj�G;?"~�՗�Ѥ�����T��b��Z��p졙&��T*7~����9�<{)�z4�1~%���a۬#�
���ً�@?� 4�\�]��xN=n<�`nO%� �_A�ĥ#-ei��--�05v�|���`�]Kg�	��Ծ��#���H����\��$9�Пj��]{�@�;������0�S_���SG��]�Plɖ`{��TmTǫ e,����45{�����	�N&F_�׬]H�V�p�cW��M�*�4����͌zw/��25IL�9[�%C(�����Ԟ"mq\�����r��}HPLG>���D&ѥ�W|��l�|�,���8v�|K9��HН(%�4ߵ �,���܇�����cպ�D�B�
�Q��U8YG���]�U�ʂ��{��$�Q+�+ŴP��ߡ1c\hiu�^��s_u���y
����l> ��L��W��.4��lS�y�0�:1g�`\T�%X�L�g��u�.�H��9|uJ�Z���^�-˧�~S�!��V�0Z2<S~��c��īz��nK>XGӾ4�rCbBYZ�D|���G����֦����Q�n@!�}N�����QI�ǲL���Ռ�'v�������!��eQ[�X�̓��@Q��Ř�m����0:a���� +p�A��Drd�	!������%~���7����Sɦ�tG|��(��2� �A�ȫ�%g��|���zL)�K���#/�,���>�?��>Oӳ�]y��L�y�#�|��pM�b��O �vUͭ�p��^B���h�r�<���7tn��$V	��(Z_I$ݶ�|�����!h�l{^��l	m@W���u=��(�2un9%�Nv#k�	��I0�$�$���erD���(d鞉��k���R�sEw:j5�+�K���e�U}6aj���-��&�*�BG��fֳ{�� �V>�'@��' P�rê���%�i�v���;�0�S�,?��_�7<�}�/��0\��@���͂K�Yj3h����ݽ>�R�&v������{�T���h�p�y���H�-O#���5 �8�LP��i (��o��]�m�?�����*�."ҞăS�Dx�&q(Cm��zN�bg���Z^`��}.+~�x�jS�e6��BYIl��*љ��&��m���E:W��9�d�?t��෮.�S�h����_����[�*+���^_�j?�J�x�l�eC�O*���s�c�����7�%iv��εY����녓a��r)
Rj�#�}�ɿ� I�����AHo{����G��X�����I�uTC���L�\?~���ߑ#L+В����&��7r+���%b�Om�*�H9��O����ؚ<�0�k&�\y�Wٷ�W�Q7or7r_���a6�|�>�)iP��.��O$�S�>��P,����;�~�����H�p�'Z��6^2�8����pb#G)X� ��u�㈤�����|o<o�%����2�0�kGϲlA0j�>I1��N�v��O�:��_��0���#�PG�hRL����y�����8�hlhnZHE�1���t$�Reߓ��F8D���9