��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!��ߌn��-��,cF�W���oS�\7b��&7����p��N�u�25��D�l�W�=%�1�Q�jzk��Ŷ_��s��Ȓ��{���������
yKR��P�*��*�8-�A�)�ӪRG� �j~����:Gd.�TB��C�m���`�ʰ�l\��/-��W&�R��ѯ�OP2�>�Ƥ��Թ�?����~}=c�3K*Un����4YG/'1�B(N����Ҝ���.�ߢ��fŴWٰo��|���"�������L�l�F֍]"���zsv��D{�yt�t�{u��͏B
 9u�J���:>(P��-�[޲|Y��zkօ�1^�vC�$VH#�$������%M;����,rq��.����*��ȿ�OS8��Z�48����t��)�q��A�����e���{�c��B�%l�
���7�ƙ�c�T6�u�5�������,ѠH�K�\������l��˛qO#̻��rKjf) t��oν���I@*@���{�P�$�g�:��^8)�v�rZ���	dI�i����/��UP%%��ԋKm��{��,�{<;���4�u:[$���%<�z�Ȉ�h�)3ȯ��~�sHrK��AҨSU�m\"Q���
Z���J�%���Ρ%�s`P�yL��h�V<Lrk�B5�v��r�h+�Q(\��mJ����I9
KB�~�p#ZP�c ���|4���7ġz�v��!Z�sX�����;��!D����N���@����eJ3�}O�w�1�m��0.�]X���l��fc�/�s�d
$taFx�-���.E$���o��b���T�]���A�qU?o�z��S~��q)��i�jD4�(\��,^[����>��,���/���{���8���w���-���ǹPE�#���<��b�f�x�x369�@�[i^�F����q{�;Cm}�)z�G�@jT��=a�W���?�J��&�!(3�K,��,z1Q�i�F�0͝q�ĭ�7�i�?p��.{�h�V6Os.�����41^Q>[�� �	�[H�Fh�U�c��S��f�_+%r�L�XP"/u]�V�����K=o,���J0�|-�`��Z�;�i��e��:]�����#���;Y�A���2��%���]���Y>�
��:[S!"�٬�5����ݚ��d��	m^i!�͆��� �t�c�<!<�i-}�&No��$ʋ|�MD��,Y|��'
�*6��3ҡ��qw:Y���6T�%��ػ={f���L��
,b���d���E8�e�y2�@�Cc������ͥ�ʴ [aI?�#� �AN(���7�J[�>���	<E=?�E;.��[�Z!&���d�V"h��?�{9�5�"(r,��{/�V%+Ɏ8��3���o��d��H����\�K��	i.ǭ߅�F��M�|{����(�m�s�Lt��%�YQ� :0��#!78 a��}��"5��%
�ۉU�&���}�2�Vʤ�X�$���U�d�x�f��7	���5�06���όg�Ct�T"=�C07`I�'�A�̶�{x��ܭ�xE�e�ŋKjQ.�ƿA��R ���m�@�L g<���W�4���SM�v�|�Z1��8��p��ɔ����W����
e2+��p���!�*��d@3�^ ��Du���H�y�Y�'�8��G�k}�?`����,�ٱhVo�ǂd�]����C�|;_G�5�t~~\���G�J�8?���KT�Z`��w&��_�fM~*�q�������%Ѐ)�A��C���Z�h�/��[�'��1,�G��3|:7l�D/8_&*��J^$��P$�<(l�J(i-��.i�<�N�C!��df��I۶��X�KF.��c�B�2�o�;a��}0$%{W�M��]ޝݦS�C�p��=�ۚ��yj��H��YF�|o�Uϼ)�g�
���cON����z��:���~��|a�Z�͐Y-���^������| ��?�ͩ�B�:����L�y�R�%�Y�uQA�S4��B�u�(�ʴ�!K,����`���g}%��Ι*�Ҥ���拾���<
\����q�5�	��/�Lz��	��Y��*���	{z�x6��ԡ�{k�Ԥ���]���T�:�-6<��e��ǷF;��c���!!g����˓I)�~�������ö���yG�Ҥ�c#�љ��Pk�	 �^B�7b��po��"�@����㶅�_�mJ�A����� ���m��u�l�=�\Pb�A��Be�߼�T4��f������II��#�+i� c�`�,|A�1�3�� �m]�Ak���j�^0dd�!���)���BƋ��Ȫ"�O%h��5���K��DӾ�|>�qM�*JT	>�}���W�r}KgnsM
�+`�4� #ۆt�7����X��cn$���y}Pg*��`HW8�F����a��%��*~�m�djg����r�Ӌ�����Z�l0�g^g@�	�{��'�L`�P�����Ѓ��e�=$9F�"8W/�����N�5��
+'d(�M������=���(94�C�!@o=���h>���U$7l�O,���\bd�W?�'EY��{)?�	��rB�	p�׌�TA�n�&��K	h����,�hT�:������p�2���j�F��rIdPA���	4n��L{�}p��_��ɔ���_2[$��No�9p�@ҶB޳���H�D<b$��ZqV�B+�+�,���q����:*G�>����b/Q�vjRŘ;#� ��(���4����	ag��}Id���N�|c�Ϣ�"�{�D	N͚�_/�O�`�xA�}q�F��z��t����� ��Jq��P�<�Ӽ����r�M2KZ=�~�Ǹ`���G8��U������C�h=��uO��	��C�Qm]3e����NX��x�щF�%ت�v/v���j?0�`xQ��k�=K�/o�m���x�x�MTgF�II�쭙A-�VS,2���?�v>�B����Ǩ0cjТGP|��$~� �oZ�rzҨ��W��/)3�ς����Ś���)u$��:e^�r8!nk-ׯ4h�b�-Y�!f<Ḧ�z�T�g��\��\�c5�����IR$Ԧ�X���/p�d�>q�\�kM��"�'��Y�|~�0��s��)k����>V'��]W�D��Nt�.E��	%�|j&(h]n�{���Z��/M4L2MT��2Z���XI�Rw���Ȭ�4pgH��>����x�K�����L�d����6�.̿a�����ؤ�tc�u�� �=c��	�A��'*���C�~DS7���� ťBrT;F��0�Yqga߂���.�&GA�şc�~2� IҞ��Ί6&E���L`	ŵuu���B��@���J�s�c��M(�~��a�p (B�"2�y�X��%��]_&�s㤺�F�ְ��c��)�wbP���Ò�V�o���W���6Q���t�E��6�]3�I�J�R�巎�}��q&.��=af�O�r���p��@�pn3<�:���(��!r��f�'�BU}KJ��#*T��=���u�J�a���]�WL1��X�x�=��A[�'fWy��iI�A� Ev�[̐��7�;�C\�Īv:���h	ADfI`i¸�����q���IW$�i�Ny>�tHﶕF���S#���{.���>T�z�(ԁ��"#D�]�Pc�H2��tj���M�Ms�$��5�������6xQ�h���m�.{0��i�%&XJ��xc{�%7��(j&����`9h�]�f4��&@L ��O�̲�.��	�+A�0�/1:���Ȁ-�ڂ�O9櫍��i#�����$��[I<1_�l b��T�:;۰]��X��I��1�)�5>��+�qpn@��>|�>K!tF-%IG1}$�:sR�\�ͪ#f�Aө�
��S�#�+(�G��Y������W��ď�@b�] �9�43�#���@�'f��7��q&���4j��l�2k�e�J]���[`��ǧv.4��|8)�6&���,�ت�إL`Q���-��P��4�ڃC���h9G�
���(�Q.k8���u��J:QLj\�����C^�dq_Y�-���ƒ���z�x�\�_JL��n��#�g�|*�]T!���ϐ2�����ͦ��_�o�{,��c��H4���E�o��!|QkM�Bn�L�!�Z	�ݻFdp�I�Oi �A�~ځ�������py���ӝQ���GC���yP��FT�v�g���WGR��qm��Vy[�V4� �^+�sL�m9��)Mf0_��C�W�sM:X���۰���mQb�t_/[�S���ݦR�]ǋR�Xz��y�-��U��!-�.hrp���s�\�H�XD�gz�ͫ�;>]l\k��"�V��<�Z!�S� �U/~�/=�k�^-�.��o-�����Y'�	F�$��)qOG��z����Gt�0�+:Og�N�:hP
'V~R�ܬ�%**Vݽ[��>�*�I.b8l�l��y{��.���fM��{
�<6��<hԏW�[�Q�W���ԥ����A�l�v�j^��}Y���r��ݻF4����p��Tp�<�������̡�m��[f��?^����+�Y�k��FTL�����AQ9�����{���=b�� �	��Lk��88��.&l��r�ڝ�0��R\j��}�m�Gŝ�J�5̈́G��S�~�tt�IXs���/s�>c�"�����E���3�F��C�C2�,{��aY��v�}�I2���w�O���o��u�
�%K�d3GG�P~�5�M��~�S�}�Z�)�4�@��is�s�z�;ث��1"),�w.�%�����?X^u%EІ`2��὜>�	.�P�wT��R
�xb�8@o/��jMп��%�~q���pj�Kh�k��_ C��sdov�Xޒ�<�����{��{̬HT,�i��w:�w
	�b��8ǯT:�ὥ�na��2��z��#������E��WgP���u�/�dN���ۘ���������_7{����JQ/oA���(�&7��>=��P�Q���X���ڍݜ4�zZ�<kf��y�epAM�sj ���K3��=�mU�Ρ��ֹT�+E�a�&F�-���_~�,���s�_��</�QG���ʨbˌB�{F3n�&�ej��w��0�.+�? <�+H��Nݴ�
oWFCT��	�~09�Q��kX攟��,_��<>~m	��N_��3�Ke�}���;�*��<�J�0���nY���U��������V!��sD%6�����|��d��dm���W������Nu}r!^0I�V�SH�5��r� ��A1�e"hK�=�<�+���&p��'d<�'�����nڵm��w��FO㣭S��C��k�x$�@�;�}d���So6@bvb�~���H��-\�&���9�n���IW4��L��+�O;��W�����ӂ R��kw��?)�i��b��-�j3�R������ /��k�Ϡ��GWF������pfy�q(�kyT�Iv[bc_ZY�<��� r�6�j��䭿1�μd�to'gx@��C�ѧ&�r����]l�O�c�x'�WT.GOe������/jn����$��y����Ȯ��Yz�|��C�,e��uD;'�������E�4��oJV�$�������z\���%loA�6g;c���Zr�~ds��}��p�|�����r���.�\&���]*\�2%�9>[���C�T��Y�@-LHp<[0��KV~j��~Tn���7u�]�!箑��3q���>M�+�$}�:� WD�[�U�>m���@7�u@Q�gF��F��^_r@@�g�i�h����A$-�f�y,A�Zͣ��)�9��f�޿�]f�g#Jr�5�w�X���өd|�����,52��P�3Jڜ�u�1���~��%,�&�Bm�<lhY;Oܰaa�	��
��\M t�ib�:p|�@�T��G��*�>/IH�و�p��.]����;�/���x�)%�<����[h�7�#��ܩSIBe}IX��L�"^,�������)��bx�:�;���d+w��(�NI]���=��夋e̻X��H�����UPâ^��T�Q��D�UH�9 �B�D�~� ^�P��~G=�܎�*���4>�T���4w�es$�8������<����#{�&ay���YIe��О��E����ڙI�	Mٿ6X�d���ٚ��6���e�J9'O��UZ�#l�%�>)��&��BZ�٠ܮz��lz9a�M�e���G:9��t��X8x��}
>��D� I�}��_)SQ>�'m�<�>����A��&Fj�ߣ�з����U�Vdme��s�L� �@�C-���BZ�`��.w�?8\4Ftd�d���-�O
X�!>ҩ v�YF��LJ��6����kJ���x��s������<g5L?*�n���!$���ɳ4��k��D�)Y��������Q���A/�W��'�D8j���G2�̨z5�qElę���Aj�1HT+e�u�D)HL��aF��XZLF�Z1Z	��	���m������k�3���;LT�
5� �y��w>E8zG�w�������:�Yo?�`L��5N��Z3q/+�+-Y M2��o1&ް�EdJ0����9Fi7I=��dK���m27>�M��HL��Y�@n��&;t0�!�P�	��K:H�����j��t:y	��0U���z�(Օ{�j;�hV������X �P�que�KH�B��
�_� �HY8��\o���oٲ�.g�������eq����"�å��I1�>�B�Ͳ�2w�����>=H���@�db@P{�D䢤8��;jW�WD|�S��̔W d3BS�B�1ýfW	?cz��rܪ��c��:p$�_Й�j14M8zp�x�t/�K>�a�ig3��K�け�Oϛ��X!XU���$�Q�=�GK�����QKcX�q�BT�y�q�ee�)B&�Z�N�,v�Ɇ@	���AǡqR�����Ah�UDQ���e�[�BU6=+ڊ���`"0+�����e�.lj��r�)=��$����KB�v-M֯������2(��_�B�IY�o4�Ѫ2���^R��mq?���j�<�G,IK��H��[���Bκ�+ֻ{b�rكk1o��ҍ�L��z�*�O�UB��~�]��PBc��m�%����y(YqHj�qkY`i���Or��n;�YX��X�7\},���y�u�!���̞M~�;#Rb��������r�	6� @�#�!;Z8�\��:�Yګ��&��*��~l�|��c�F�_]�J��r��B��l��a�Z��I�uR.�j�iv�_�\�dc��E�e��+�2��J�s��\	�@8vUP�ߘK��3I!��%��E��녌����0������7ô^��*����	�Ⲅ������U�͕b��0'�8>�H����Ń���ܳ����6��
���PAa���9�BN@K����M0��{�������&a��R;	�s�b���/�����^�������zȉ#�NCSAY�6�[B�|��r�//�*^"+f7�em�>r�/����iø,�o#�X..o�B�I�U��cx}��I�����>��sX#��;�a[:&!dm^��-�z/x��q7F�;�����)]V�hB�Gi�v��$?��۫�[�Ҍ�Z�����\ݢ�l�Dd�7S��:�v���9������#��~*��r����rQ��5N,�JaTޡ����*��	{�G�ĤT��|�D���@�j>%P��$g��VZ�l$C�7b��9q �����e�B�V�6sM�гt�csK0����} N@گO���cHWO[����V爰�s��,�^0L�\��Uv��m�UE~�䣒\�B�l�Y6��Ŵ��mw�(]��3���Q�)|��gcJ	�g�gz��[u:қ>Y�A��	�ip^��Ʉ.%�nl��3	G%h����"�U��r�zs$��7������J
��72���r(s'��W��p�{d>MPF`�T�E޻@��z���]��~+k��n��DK�U1�'1��,�)d!|Im���t�+�����Е�<�N ��b<�jI Tsf�/ ډ"��.!~�~�4Qvx�+���A h���=�x_Z�mŇ�����o�F��ep����i?��<v�w �r���V�d��]���+��n���|w�6`���n:3�� ov�#���B�	����-5�ֵ!O�g1��\N��$c`,j�W9���:$Ĕ}���荘(�;�_�M���/�G&u'_��1z4��3�O�cd��ĩ~ި�'��0���>�ˣ$`��C���3<�M�� �e�rЀ�2�.�bq�r��W�ZF<9�_�R1�����I��~��EB�O(!^8��ܵk�p�M[6�ת󣊣i�UT�MJ���	�C�u��lS%+'Q�'E����6�DLjJ�󿆲.��<[�I��2nPv�<w�ٯCk����?�S�k�.�)�c����B�1 �E� �ԥ
�ؘ X��m���>$ᕠ".ݳ�11�_ٟڇV�HJ��#L��%�e�����u&9~���y�s�/�h��ǬB[���p�5\7��ф��<�\Q�� �L��<ѐΙ��h۳��@]a�b�N �n]�z޼	>��I�;6�p��C���[���b{�6�w$�K�}v��f��tҶ�����&�B�z4�V�]v����.��8ҶN�o�lk�̵d�Ψ��"f|��]s�p�w�XCO�S��1����}DO{�i�E������זjh�Yh����>iu�Kpn�G���i���W��72����u�@�s_׀8~�b��Yԅ���ꭏ�"3Kߗ���̼6�[
���9�-��n�'v��H^?/L&����]0颵�*+��L���N��e��HG�Z@�x�@�3pD�����	�r�^zua��cTKՇ�#x�)�5�/�Lwg���Xtn�9�"�9��4�{/�Qv�/�J5�N���بr-�u��-(<@�ut��+ؐ����6�y���j���G�������ÉBlݛZԙ���u��>p�N�m)=��%�: B�"�q�m��)0�.�:ؽ�EP!=�Cp�/�i�/�'��1��~ ,�Q� Ə�� R����r�§]��P������h9&ģ��ӡ��7��b����o�:l�z���>3��\�T�S��,�px�����ؽ����33Q�36gO��Ɍ��aϴ��f�D�1VSت�烟Te�ȒmQNF�&�	d%J���7oڢ���Isx�^dS�w/<(v�*���J��4��b���E�?g씋�E6>Ms�x)L�Z����H�n'�x�f�:t���}�@���yL�\������j���M��ޣ�����uG�J�pD����Ｙ��~a���pB><?��! �S(4��o��h��}��;��S=�� s h�ɕ�Ϳ���O��U���)�:'��7��o�p-���R��\S�s��h���342�wm�@��� ��MA>��X�=��`���Y娄d#y��D��1��g�	(�<ϑ����$£�Pz�	&*�M��j�Ge5���x򅅹��k7�pZ�S���?�Jk������ RA1F��H�=)�qc�0]&�x�kR-l@�
3�
�ǟ��� /@��E.ԩQb\KM��1���i�pF0��ނ|/S������+�t����_�=ٿ�ӑ�����0��/����5�4����%����2Z�٩p��ȸ|�7�e��AOe������ϛp�&��Aᷜ�xBY|�E%@�^��L�GZ?��yѫ�o��Ŋ�.Q���>aՁ�J89�� ���c[���5��ȶ_�b�x��cW3�O�D{�vs��^w)"�e����o4��l��ט+,X;v2da㒨�&]wt����|��7K�K� d���J  �B=����q!�kl�#�Z-BBb��7�dS����Ǯ��c|�����m�PW��U�T�A�s�Yh��j�5{�N����d��@��D�o$>vC�;EK�\-㰑�|���a����UW�pa�fL������e�:�T�:/�~Q͜p�"y�5�<ȝ�Ԏ���{�u�*��o��q����Q����3HZY���߿i��m 0:�8L~��]���t�}�hyث��*�4�<�h�Ɂ0J�[т�>����/��)�M�v��#G����������ԗaXR����B�&�90�����b���뭇PS��4���9o��j>y�"+=-\L��&�&a��kc�D�u�Syd�鰲��E:>��&�7���[�o�9��n�P��ۨ��O�"�?�W�@Q�8Ֆڥ^���F���1͝|ꬨat�D�hA���v9�s�<�:��a�
�B�1ݻ�J����L���M�q�Y�LO�'ͩu<85;�^�Sm��TN��K,c�1�2�f���:���$q?6�I��I`X�����Wi�Hs���$"�����w�:u4Mr�@��l�"=s���S[�>{$P���U����ǉ��c��I3�Đ����*�"��g8]�d��6X���V�s,ܞC.R����7\����3+	�����rG�*�,99�2��ڦ�FZH��	1^y�RӰ�;�H�����Đ�F�|b�������5F����U���� W����`ױ����F�Cm�0K�}�s����,����/