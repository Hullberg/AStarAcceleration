��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!��ߌ�6�u��S�`T
��E�E� -�5x8�ym�7�4�����Ƹ˲[�B�?�O�a4�����ȅ~��>����8.�NSTiӸ-s�M��(��1��4{Bm}j�o��#�,�.F`�_S製H����;�!w|] ��{/IK�����_�k�h�Ci/qS�� +P|,��WX;89zq1��f[���_���뷭��`n� �i.pW���Hog��/a�pD��+�;k��K@5�����5�O�XR#����J�9���Jz-J-��B�1��gI�N���I��	�M-E])W+ 4~-�]��T�vQ>C��c!°S�+MjB��s�#�N�˔#��xT�jQ�ʀ�q]6�C����Y^��*�<���IpP���C���&"�C���c��_M"����� b��v����4xe	��	p����B �*=I�j�E����x󌒮�b���ڙq��hQ��$�}�z,�ϩ� �G
����R4����:Kr�-��qx��N��S�'��t�=[+�rb��#�xt�H��T8
���Q�	~���V�Of����N��E<LiZ��a��n`�����~���ҟв��bѺ)�V��B���$�ǓRnN+{����5�Q��$R���Z �^-� 9I�LN����	��?����B����_\�XF+�[G�"��@
d�;VQ�F���w�O(���co�b��-{�}�u��7J1��%�n���?�ex�K�K�`C�"IK�Jg�}"tRc�$"�J�� F:j��8T�mD?�G�!X�=�Ρ*w�N��A�lm��h��J��|B��'�
�'�CM���E�l�>�UK����4��a=.�*�BP����+���ӿ2��֜�޷����]v��M�a�am� N0�l�;.bO`�/k��C�vY�E~�d��4J����t��eZ�)�@�M��$���p��-n��Ph��^�/���hn4M����Y z9�=���� W.~"��cUcm�ߒ��`�Fg�=F���Z_];��	�PsƊ^���=ǩe@	q����8��h3YU��\]I*�Hؙ̻����|��4$ �` KCq��w+�g�����jâ�>	j��f� T'7���6�_��Kּ9q��b��v�.@�5�]���9�U�h�Ϻ=%���6RK�S\���G���F��v��fڔs
�_�U�J�����pdβ��uUS��~�d�]�U=!Y��~�g��|�ֿ���_�ͷ'����<���&�s��@'`�;��0%�>�ro�r`���?u��m3���hL����TMP�Y�K\��o�R�R��4��(��e�}��� ���;H>���Η01���'?_k�K(�Dy�����t�̔b.����v4O�v�b�VԱ5���[����62��Ԏ;��U~t��Cg����+��zK��z�^��ƞ��t���̊\�'��k�?�"$'o q�K���5�pK;s���|�j�B{�	z.2�&Ҭ��&�g,O�oor���dLI����H���!�H�[���4��u�v�2r�V����yvu�?M�P87����]A�B��濌�uIο�J��z;�*_�X�~�̝e��9N9A��ȴ0�:��_���À��K��BP���F��A���`�u��J��<m�~i�����|z��%�ļ	1��e#����s���6�[*���zN (�L������&cO�ph�V�Ny�[җ������W%��� T����B@�qh�f7��d!7�ع�>d�������c����JQ��fKy�������N�b�a1Ctx�Ofw���凮C���n�(�?8��6�c�/���J�Ր�ښ ظ9
	 ������>nO<(�P��[��  �����k�֖d��N	'ي��n�M���°+yfs}*�]I]�Lȫ�X�S�&�zߵ��$�8�ݤN��B��!4�E��@-i{oBZ۔�j����}x(��ȷ�n*x�i�ۆ(�Int��՞J�k+��v���x+���E��%-�f}ʭ���Ќ.�q�e���yQάI�9P^�:�c	|���4����Ŭa��XۿE���0�bFd�����C����Lkg�e�{��I�l�{�mDxʸ�#WQ��,u�� ���H>��=pO4뭋Hg�F�����OO��%/���z2���V�HCt ��8s�bC�}=�[�#p>�q�0e��;O�!L�V�X�Y �;t�2F;d�-���!��[�V�h��}&^�t��ǆ�h�7'��7�f���C�3������=��/��b�A��h�1o<�8Kq�Dt�#*ԋ�����V�n�M�!;l{�	�X7�2N��	H���ӽ�F�+E���i�>�[�9��4~K�N
�.�T�Qx����Fww!���C{O�A5�q�C��Si�IV4V�#OŞ2�S2�@��g�=�P`��N��#x��x�K3�-��'�,y`F6��B� ޮ��%w>)R�.5Ac8y�쟨��!JAT�m�&u*k��o��e%G��4q
$�W�Ɉq!���n*��K��du�0���C:,�' �}��q��|�!��U *�?g�Ib�t�p%��~�|�ZH��=zTGs��Q$x������(�����	�m" �����Iu��l�p`ƣ8��h;
������>z�6�f�hņt���>��;�e�w�aj�'�yL���,�Io,}�[H�S�R<n�{u_�����7	x�%RR�L<Dd��T�7I�~��e����Z�s�d{{�X��	H
E��|wXd
i�B�T��/3;�����M���#����V80B��a����F����)�����N%�>�JGz��?),�q�cO8�@��Ӭ�K�[Y���vT!�T<3����4�x+��5�K�	�)x��?�ڂّ��>t�<�՝���CBcN�:ʉUU����o��$����� w
�x e��V��&�o9-��RU�S����_�Bf�c�ޅ�.B��Z�Kq;�e@��M�Bo�����4�H4���/�M����Z8�f�	+���If��#f�����\��Jy6�1��8Im�>�̔��7���Ld^ѓ�&����������ܨ��Z�9����(QR��3��B��l�9mK�27g���5ׂ���܁Z譴�
E���+����$��Cd1��CL &��^�2lE�]5rN��ZQP��T�P�����)i�W��ґ#��d�`S0���v��%ai��(˴w	��*]�$�4Z�Œ"�1��y"$SLMR�i��cr�P���&k2�9 �8�l�������"�̓h"��N�P[V(�&I߂�>�qҴ��GS"r����.G;T��O�|rU��$Ŷb��)�;Z�]�;��e���`d��u#�����wZ�5�݉2��C6��"S~��U���,��:�1��sB���X�S�$(cW�YaC�}�F�~�������l�)q�S�@����x��L���B~�}�#�2���oR��Et^rL���-�����-&,j�����`'	>�Y�+Q�}�([� ;*�3m�&���Sގ� ��Ӆ�5;����b����R�w�� ��S[K�t��³��$�"ǃqDg�fKQ7WO�E��2��G������O[{��~�V1hA"+Rl�]�JF�.�.~���p���'�$�?�Fo7k�u6	p��rm�SC���;؍��sBI2��l$�&��b��rŇP�$�'��� d@����V��P���~G�e�;�,�B��v�����ū����zF]`"w[��{d/�:*ڔ�B��T��|LiU�o3�����aE3�@E �RM[�H]�Vr W��lI�;g��"��̀%�1]���7o�m�l�N��=��m���k��_�������*hӄ���}��q��E�i���'m�i�_l�3pǡ�O�d#��ML�xB~�	ٞ ]��֫�MR[�
�6��;sI��|��.}/]�׮�	����+;kC4�pj�}��kjR�����I��0(\y�8?�`�s�ʑ�Lyxo]b����Ee�w꽪��
�qQ�Nޖ¼���aѵE�:�Z0g�L�#>+��!�Zk��v���(�	:t�h��P�"[8��䘄���xu��>
Z��w��_���U�H�=0����� -g�/T�;��}��s��O��YI���P	��Ԟ�=���C(y���ڋá6C��K�=ό;�J(�1��`a��ɜx�Yp�����8;�o[9t��w�9ĳ(ܦ����XU���=bo�}��ЯIYG�S���@F��+є;'��>����Ef
)��	�!d[�4-56q�	���E�'=g�Q���v#e�a<E�䉛N�����;�� * �'��1�&_܍h@�ٴa�V4�ABUlC���KM���l��l���VF���������7�H+��`8�ZPd�Ѩ�j�C��甩�#�:�1��"��1r�{�i!�&VP3��������#1*��a^�Z2r����1�$Sye����G�]�j�"�G�
/�!6V�%G��^�=���r��xC!�j����b�� a��3*R�: �b8�5����ѩx�Z��ٜ�2:J�O�%lb��@V�����\I�^�>�9���VP�BM�S#������!\Y/���)�Sԝ�78�W�lh�aRU{ќ��g�s��L�8r�<cu=��P�j�0ȭ�q��N�"o	t� �Z�m)y�	q3E�1RK����]�[3�v�w�;�?��m�vzЂ��\x�l�!�v��UC� ��4My4C#��6��ݞE�.i��̇�Q�a^g��8�ƒ�}���8,�_S��49���b�Ծ`gz
�
~H�d��ݖ}�%��T�4͘����vW��S�ϴդ��t/��j�ˁj,\QZ��XMX���K�!(��bɹ�t1��.3T���ӭm%?��NZ��*�fQ�<���ѣ�����A0��z�w_�t׀/A{7�K�C׏cZ�	Dk@b���A�B���}�3��"�K5��`�6*i�(��/�����j�3��]O��`�p��
D���<.��~�v�`������f�{�c}u��b��JヷҊua�}Ƒ�+�/2��Z����\����k��M�,^~��|JƎ-6�{q�O���߱PPv��y�S�rr����K.��	Қih��C�D�JG�
虱L!�U�����2�d˸����E� M�]�VL��v��Tf�/Ԟ�+B�
r&_�p�6E~uN�)6v�}��g�=��B��"'��Zn(�<�զw�������~W�,3_��]AC���~������]hݎ�3�K+��{�zs�*�)E��5�s�%� ��<��vMb�����N��T��}	G�|{v�c�\�� YHl�#���Ă.�
=k��v/�
�����2jsXg����h���t�#�$V�]ck���l��n���I��R*])�i�P��V;(�	jʷޡ �վ�OE�+)jLi�k:��IKp�3������:a;�1���h���2�G-p4iB@��	b}w�ι�b�W�l��������Ȃ*(�L��Z�������y���0w	��'�=���f��r���[QpA��"2�����JV����o��X��"�0��H�%w��ǽX�C�$!z���$"l�W��V��K�*`l��U�[�a������Jmb�����ε}�#�bW'�f���L��Xv�<��a��<�����>�5�`�����̂+nW�t4g�K�O�ڟ#����	 ���&��R�k��ي�'�K�k

K��ժ�ón6>ƿ�+|t��Cu��dI��)wr�{<"��e��g�c_��QtVl� ��v!�
VWgsiY���L��㮾'��t]g�c���K=5�^�5�"9��]�O��!s9��"��:�)O�e��jN�)sw��Bڊ��U);�8
�iZqR�q���e=���Bp� ~>�PL���7�u��Y�O�
�1��Gb*?)��0f�p��_�����ڴ�N�/\x���"Fl�h�����
���Z��w�OQ��^�h�����b��V�@S�U��|�ʺ�g�r�t�#6��}��ɸ����DV�*ː��G�0g����.A:�1�W"���Ð�%�;�y>��u���)�2MD@>�+�$�M,�����s��Ǻ,v��� �9��jʮ|��r��S�꣏�F�00�ϻ��Xt�rt��J
<��7���E�����=�iÆwv�q�j�#k*��%�k"x�k�����gGPVe�7r�珬`��t0_cx�&Ù���z����~ۨ5t@`�}���dG�_��T@^����8���@�m��f��É����42��Ğ!>�3a�q
�<�G�� HI�co{y�Y;i��o�a��ԹȆQ(D��H�%��Dv�M�Y!����&��!�4�ꔹ�F���Z�-��w����������iq���S�g�E.U���֓�����T{ZheE$ȵ[ƑKH͂�h��tƵ:
K��ުk]��I���E�~W�VJ�MhxW��Բ}c����I�ݒq��$��t=Ģ�O7KyY�QD�TF�f��l��[����+
�	2�ڱ�bn~��t�z�!�ҟ�R4��5T[Z�)}�MbM9��r��/$�q !��p�ڕf��K���˳�#�;M��D��x��¬�]�@E���rO.~s�o%߇���Z�N�y���1K�5����z���3����W[��G'��Uc����Yd��h{ŕK0Ts[x���1��G�n�\C�����wF�W�AQ9�չ��д=������x��?�h���v����!<0BQ^*���:�'Gb��Ep���;�yKˇA��I^��b��*�h��'�j�10<�������e�K� ��g�.h������0���S�{�餴��4��CU�.�_�jՠ����FgG�͉��u-�o�x�kLc�	x� �w���*Q^�+��l��f�5�]~A?���G����;�����X.T����TE���<�4:UT�ƭ-L3H�m�� a�Exy�������翳<�bq+'��R�!��c�4��[Yt��`�*)��g~��Y��>��������,"���L��.'�t���p�!�%-�h����ؽ���,v��5���=��*\x� ��T��:xXL�{C�����d��Fe��$i��p^�5\�[x�~�&P�Hs�2��?L#�j%"N.W^B�jU��tU?�u��>	��g9��V�.3ɺWu�]4~ɫР�R��%c�+��x;��v������s�7�Q+�J�wj�s��;�W�o~�D���#��%Y6��>�4���I���g/�ׁӽ���8/��V�6M��*줴�,`\=N/��V
w~������/ӑ=��l.O�S��L(
Ŵr_l��s��>�-�S�Gy� ��;ҷ��*6}u ���g֔��{���-u	l�r�z<*�|~0y��y����97dG]C�mb��5[��F�����M��p+�	�ȶ�;��6>?�I��F�u��5�XY��x�ĝ�f��p}ߚ���J�����C-�"����W|5|q|3.$�N��5Zs�4@}�f䁽�y��Dތ�w�Y���=O��Y��l����KP]���ao���@
`�c��Qг���A�Z2յ���R؏�զg4B��JհO_����h&���Z�𚹥ެ���S?�P�g�/˯�$su���1��<����<)��ӡI��S�5����W/���glc����� ���Xj�H�������o�M7 �� a]�&H���Ge�i.W�%X�-_��n�CqZh�oݑ��M���q�c��IX�M1�^NP�toj�i(Nk3�Ŕc%�k�Z�l�/e(ZQECJD9�T��4����yiI��o4����5���Y$pf��7��k�.�����k9R�Y�mȧ���'���o�-S�8��W��jsQ�K6�*?�Zy�n?锄��^a�
�3L�D"9��)�Гw)��e�F ��B�ðY	���\��{64m>�@�`�a��h`�8�E�&ei9�Е��`)
��@�u)'C�ꉽf�X>$OY�q�/�$����IIX��M��q���-���U��6ɠ\�ߨc(�D��^�x��=Ⱥ��PSR�ǉ���3�C��
vˎ�_� �k�Q���(�9�Ñ����Czj��rN�ȾjsN{N͚�ӥ��O�����	�W|K�u1���M;$���R�9���/�{�{AV��ս�]z�-_y3p�d�nh粋�����S�oI�ل)�붏L��U�y2�������UHnqt[���� /�R��;w�!;�!R+��R�<灟�2��:ÂV�,����ГS��%og��J3Zs�e��n��i&՘0��:�Fkk{��u.pu������ݜcE��eo64�}�;n���(]a%�gc ��Eօ`S��Dw��g@b��Lgfbv�"c �s�5�*栚�7Uҝ�������)�)�ƌ�NŇ�.�ow�y>C�_���z�<��S�ܭk��w����Z�x1�@-�E���
ܾn�����_�sP�(uM���B}�����	[5���'�7�,5��r��}��T�8�>Ԑpz6��x���A���5�fXj����a�71���b�B<����%��ͫ�����%�蓒$���M�K��_J���nN�0rrT�]��KM�t���LDc�V�":m�xQ�����>���,}7W֖�F�C�d��Ӣ��p���V�#���,��J{5i�3�\� g4��⩆�EV��+��TZ�*�F`�������TM��/�b�$bO��u�	���N�ͻ�H������%�:��hU=��	�rV�>2��ڳ�p��;of�ʽD�J�!��Yfњh��7Y���xl����Ţ�|m��񻸠_�H�4t��Z�2! M��"n^������x�%��LF���<�Q���u}} ��Z#W՞^=�JDh�s1L���jDЍ}����jP9ѿ�^��8��*��,a�Zg�Ť�s��8^�ɰ2P�p��iv"yC�-
��kIKS��E�FD�*-���c�>�i�G�N׶���9�n�