��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸�Σ�HڂͨgT�W�1�.�gW(�CpzQx�E�.^F�tZ�����t�I�k+ǉ������]�+����a�5�����^���b`�	9G�2�Pڵ�)�K5Xi���o�	վW31؁�����N?���r{����M���m�(p�׎!_�:�f������K�q�)`u�E�u50��� �,6>���76w޻����3�����o�ɿs��@ܤ�ۿ�fц����=U/AJ�Y�z7KKG�S6�PniJa��z�k�¾;%�O�Dx|�e����,�Z���}��:��X?�l���Mr�b���'|-��7��s̊.�wiQ�__2�l2��C�.i�7~�YM��ؼ�wJ���> �uB]�>1sR��w2�Q ����~VM��౦�Zp�8 h F�����J$�P:cʕ�t�.xmyr����8yg�"�����lF_ �����+�b�J�� Q���l�T�j)��/d�ϼo�p�w����"i즌ݺv�� qk���ިxڮ}JIb1�}Ϲ��9䫽�kO��VlD֝��Ӫ�P����O�^��$Y�]$}3ʊfv��!W��F6k`�!nb�S�&hE��$��ob�g�t�5��F��/ ~����]ƭ�&�~��s�ź� ��[Tl�H�w��X/��N+nz�2�X�`C�Z���?"@6-s�F��j5��q��}�/'�z�ٍ�Eӝ�o˯4�,�7��];9��Q%��Bz�zN���`S�f(�m��m����"E����¿ڗL%�MJ��Q:��JR�L���QrR�;�-��;���>>�d�]����qƊU�}�E''��}" ���tg�wG�%�=��{�	a�6Ǡ��ɪ�H�b�~���WEzͿۛP�@��Im��Ε�=][�|g�Z�n��e���۝
�Az!�Z=a��%Љ��=�Eއ^�HƫLXĆʜy�6d�����g4�e��Zё[g©dQؑ��{z�z��6vZ��:0UP�e�%00�Y�+5+=1iH�F��h��?�@��J;{��w0�ʘ�WD�;q&��dG#��퇨��Ж4L�|����u5�q&�Q�����2Y��cg�DG7
t�tE��|��z�3�J*��O��?YN��3h�<��ť��l��Ju��9�F��!�G&��%Ǚx	$	��hVl�=�Fvu{&�O��!"�y�u֢:�"��ȑ�E|� �s�Z�l_Q��\d�|/����Z���l»�O����5�%B�J��:(sdF���ƺ��ۭ-p[�ZQ+<(�n�Pw]NB:ۥvn�*�"2CR�-�N+5#�_��>���4f+�$��^�q�X����\��(ɿ�X�
_���a�]��_��㕞/qw����I]��"�s�πX(���ѐ��SYןƐ	|����Df���_�,ݓ�i9I�u>��s�{1��U���~̀h=��<��J�6�t˾���S�xI�[ן�O+Q����銱�+�岬�5L�^��}����V@�����*�i�<����D�4��+f�������s�80��Ւn/a��7�����*l���iً��r��8��;l�h`*R"����Bg%X��'t2k��`�ґ�]��x����W��z�+X5銮+��"/�EGMn�t��_��򺁂����τ������qﬄ�A4���/�xĭO�2*ﬤ0�ܧ�Q�cI�a��Ӗ��h|m"�|Le���x�*��|1�Z�J�Z���X���J?�T