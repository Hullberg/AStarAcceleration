��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!���_Tr	�ĩk�P3�W�W!���22�m�@9'X.A���������Wq�U9D�qKn�0����L@�?�ɝ�
	��$L�����4t�n��!��[����ÞJr�[@�(Q� ٔJB���sB��X
�<�=p@�<���n��d�q�����Z���)��fi�� �7y
T̚�� �|0�Ьd|�=q̯�a�.��е�%�c,�*�x��Qm���\��N�i�؁T�*�tV�m�Xd1y�	\0ŵlAw���D�
��0}�P�T��_jmP���b�J�k�!���JƘ[�D���84w8��w�����mPV�x���qX=ƛ{��FƩ�>K=��9`��l��R��yY�������������e���1􆘂�W���[r6m�3�o�0�
@1,�&�����8x��S��mP��TS� � ��^/���g2 å���d�6��"�}Gs��ENE�A �>�	ݴ�e��q�|������e�S���˦ ��ں����Ё����-c�z�a�����P�l���s��N{�Sp�J¿���sF�q ����s	}\��%W���O��ƨ�+��أV�Y�>�3T��M3�\LS��@^�9���g��l
rpF�{�5��/�&��'V�^���):�� -.?*���a���{��,�:u�^B��%��oVq�}C	��B��y�k��s~��ta�,���ݯ�/Hi|��X�k���
�cȲ*�C��X��@��绉r�	��kp���_箙���Ȃ�5b�m��8����S
������P7kG��Ma-,��5�2��^�e�.���/��ߞ�-�g_����L'�pR30�M��s����ҋ��(���$[��s�Ec���[��4&kb2�Hq9H�����R��E>6y<�ʬFJ�ڔ�S�jr�*���#�O�Y!��	5�� �����7�74꠺Ԏ�����N��"���C����כ��ZQ2GJ��f}��)�l����8>h������P�@gF�.����im��?�ʩ&|}p�@ �+)fŗB7Bt�Ԃ��s�6@��������Q�ʀ�<���E�����le����4W��`j��rȺ��I:�>��'��:�JU�*o����iFKj�x��b�%���N�1���[�&����R�&n\�jw9nR��_���}L?�|Hs�g�	�@�U�Ƽ.��&�s��1a?Rb�ZW��R=�KC��j����]JKe�m�'v��lk�hqT�����t�+�N�Ǹ�o�i&�̥U� ���H�a����[�昬G�sn�9&l�s��*�#���)��h4�}����E�\s�)��=Vk"��)P�i��Y|���T���<��P�b����pA)�{�\� �6�	�=�3��87p�U#P+G�u�u 
SV?�=��]Ry�`B��?��u?P�jP)��?��2��@W�&�X�>s�Q�]Z����@�,P9J��E,&x���P���uC�+6VR���?C(���p�2���|]U&�\
:sp�����d���_~Rł�^�����^Ϸ��7�tl�����9�f����8~��w����7��  �}Ua��.�ڧ*kR�o�N�'���2x16ɌX|n�D��y�?�g���b5K2E�\ȩ���R�@��)A�lK��׾]�YN)�4 �֡o�X)�ƾk���-�Bd��`�=�8{�v٥F����Q�֟�����_����Pyha����'2y]��݋m�P��`��ˑ�ͨ8�]v:�3__l� �?(���d�Y�	S!�պ��5�]a����6���H�"濹�����@ʾ�~v/⚴�<�3D^�����o�4)9��'�����^���f�ښ��~���pJ��gt��j��D+Ń8��f�5/����ȱ��\�q	:��R|`ɥHw��'&���K+�5o[�E�XL�	mt�ʢ�'���p0��zU��}o5�U�{݆�������2(�0w�?�C~���p!��]��������F�妯�C��7C��Fo�R�Bt��2��e�躨ĸ���m,^��p�/�k��/����HBm�j�Lvަ���1c��!��)7�z��B��um�/�W�h��'�t?���$�U{%#��D���ܰ�GW-��W��nK:������YH�g�3{[.s�����E��B��q��f ��FYB2��L�nt��S�6���=ӊ�v�7S/MMDу'���挏�������,2f4@��1�,�<�)��=懗��J�:��T�fm/�P&���E=�TA��/��
	���ּu ����/��B����%��z��
7~i�Vr���zXjd������,b{u8��ś_M����j�!�Z8頻�8� {�5�r�+׳�L�vq�8";�^\��|k]�#?�By�8�F�'