��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����
�MGZ����򏷢��+G��9R�(�q��7)�E~�3�r�c���<�)L�@$-_�\Ҹ�eM��i�2g��|7� ��,x��.N���`8����z�їM�n;
f����oEÞ|�!&M��_�U#P"u�v�����]���>d4���ƭ>�-8�֞4��h��<5[Z��|�}���ʢʜ��V%}�x�wصB,N���dT���{�4���|�����ICA#��5$)�����o�kL�h�B�1�� ��E9 �rn������ba�gR����1:0T�.�k܍�=7{#�
����dI�*�?��3�B�+D�q���ޑ��ve��F�M�w?r����_:�j�F��y��wb|Z������'t�j�&L�	�];������K��������#��b��=���əqC��d	���][[��zc�GT7��"g�N�([Ye4��[6����Rhwp��.�J����R�`2l�ܘN2��͔B�f�����]\?�M}�N(t���RG!o��!���E��lr�1���OJ��%��D)��l��٘Q놽���	􂾆*T���%�V,35����,�<
�0\́yaW�q1��
<�c����u7�3'W���S���<uށ�d[�����Ë����P"b-�{@�aX����YT����IO\f�U7,��㘌�f������{ţ����&;�B�kx� �9�����r�$���ޒg樎M���d	�DX���� ��~ze}��?O�>������p�kB
9������<�aa,P�uF�gR�,.��,uvi����~�S�0�Sd��J���R�^�6�L�7��ot�}XZo$���>|l�$J�~
�����W_N��I��.�҅�"�a5\]�$���ϫ߾{a��j{��(��EDd]�^���"���x5�F���b�V�"6�RQ�3Ԓ��+=Df[���(}�K��?�z`����(�\׍)��D�,�����)"CBq���A��ɤXP�w��9R���j�8�L�nj|r��%fN�_k�+TY�yo�	�|B�<m1�wh03Q'�d�pe0>����=����}W��d�$�5�G�L�W�Y
������1�g�Η�W��IF�8�k�_����+�
�=����f�n:2���N��އ?uT��y�_9k����ϑDm��*��Y:-s��y��=�7��_��.R~I,��8�Hj
|_��2f�ޣX���ڲ�v�>���N���
��y~{{�^AR2\�.�����i؟�s&ٕY�������'����c,}��Z��ax�A��:���.�л��̞����~����}�(��>�\��_4|����d��p�unNR��Mm�d��h*������,�u
7��������U:��H���kZ[��3V�P�	���h��:sӭ��m�E��w�G@:��>������Y�����zd){O�<��!�6��Bh�C�����=hW:L� ��<R���b���V���<��L�!�~$l.Z�`��Űi��f%��ݦ���:�;d1`���_2��LK�^	µ��ؾ?���7���i�	Aff�_t�9��Q�Ȏ-��i:Tc���"Ƽ�'���ZF�{ݍ��oUw��voh�4fЅ[yn���\�_�\�J@�2��N �J�W����$��ͣ����r5�h�ca�����w~�wE{��0��+�?�{��2��'����/�b���Yw>��� ������H��;��$k+�C�x��@>��0��)���͋�=!��>��]o��#�vh�6�-.��[�֓W�i� ������E+�	͙"$ݯ۵
.&��\���ISϬ#�J���9��7����ec�n�쒜~�]K���e"�D�D�^�[�U�1f��O�NƝL��+����+��C�!���8Pܐ�+�%���'
F�)���囹m�j�nH��tmA�S�D���#ͦ�b�?�zC��ӥ�Z.�����fB �/A��C˷s�'�B�����)�>绿�q���U �ULU�9�ErHe� ��*� .T���N����o�6��"����ؔ��j�p\���z pꭩn
�+�����g�@�q�P
�n�/�K��Z��{�6a�2r�kTn�$I��m8��Kt=�#?�7&�'��_7�s��}��#_���)��NR]9�^H��?�5�0#��4��8�;o|���$xc�h�p-�K�j�)N,��?X1Y\g�7:$�N4o���~w���%f����Q2��
�F�,�ά�����&)|I��Q���1��e#��h��j��Ry���t���Tm���C8q/F��8�4���픷Is:ó�(;i�s8�֓�pU��Ћ�ݛG���Ԗ&;��;MP�ŭ�B�Ե~%��5��ZEE�w[�����k�8��� �~�2F���Ô{��ѹp�ߙ5��7��k � p�ߌ�`9XV� I�ӓ�� o��\dw����H�T<$q@
7L��j�@L��$ϖ�^}��Xlxnǃ!�}�-JV�~�$�쥾�w�s���t�t���s�J����pܰ��?0���W/�Xo�|F[����h@��f�J�mM��6���5�7�J�NX�&<�u�~�C���I A�M�-"��@��}�.{ڞ�! Q���Cs5��d���9[]�0n��\��|l����`Ɂ��*��F��9P�������C���)��k�!~^O�״�PT���ϰkY�=]�#��<�r�Uh�M��J��qL}�h��۷�/�|Ġ�1k��~Lo'3�s��z:�O}��R�����ͼ|��{R��UӲ�0�yy�Nj��:^\"Z�������%0��0e���ME�Q9
t5(��Df�I�"�1��� ;c�R_}���D=�8����`��1q�sZ����p�sZ��`l.�w�Ab-s�V��
�V}�.��~�VG��1TAC��Ŀ8���v�R��a���0@�k�lX������W�o�8�t.ˁ���/D*&�����#�yL�&91،�t��=��C�CU�0���T��%�|bH
�1��hv<���2%�/���?㓵o=:�O�����$a���gn�����($.�{���H/�Y#cu߿�S�B���h�+���zkLb�O�s�*@�J	��%���|�����'�S�mUۜ���h�b� TlE^m/q�i$��c�������BY�����]>�rK:��cǠ��d��v-���Tʐye �؃��YA���������gV��i�s3��W�SXө�⟪��ٌ�c����w�r����J3D����$��'j ��)~��]��%	bz5ʒ�du�ɉT�K�F$^��Ӹ�+��T!1�	����};"'�MG��l�4�＋}��*XL��4�������W�F�g�f����@W��w�Y.OS���Ӗ[a����:�=�p+?]}�P�/C�S�v_�%����&�FuQ�\�Xl+���n�q����~�� �v�^�/ !-��5��\wb*���E�$_U��Q}"�\�Ї�ȇ�=�Ʀ�IpwE��Y��{}_ۃ/^*+�����d�h2��l��?ocT���e!���Vtɜ��JI����	�]���o���xg�	V�q�׬D�t�D��{�����F"�C?���"/�O_���� ��mz�	�|�����{񖇩�[T�ڃ+�@{i]�>��G��:!�!K�p����4�9�pyeV�I�T��Iw�ħ]��* ���<��V2%\<]�	h�6L����O��R]�F���/N]Ϝ`���V�=6�j:�����ÉB�5�bl���:M���=H��H͊���Kk X�(�Gq�q��A�̯�
�]��(����1��4��,{�O���ڏ�E��}0ӹ�=vLB6!W�k�YU�t]����ֶ��|L��bg��ˏ|��$f
ۙ�%�CqG�r�^|�F����@�7���U�6����rv�+�+�M��Q�DY|�$�U@g"��с�1�\��(��4�Xu�Q����S��d�h�����i0b�H+~]4�M�{#ә�$�1�;p�+\P�2��翌�Wm�^�<&��<�0�a[�__G��w�л=Y���|�̆	i�0����+H������*/=v�= ^�ȿOG���f�W�#�N��չ.��R�p	�\}K Y<5���i���Z�Ʉ� ,�;��v��Qzv��_�t��r8�N;�|	w���}��>F�j���1�j1�R��qY�~�Ĥ�g�L�E���o�QN�8�Kkư�4S��4�FC{�|�ϺY�`�D��Z� �*O�GD�^���tꀮ�K����!���]����I���2�`�]OG�%�?\�:�y��m(��ȥ
���E���x
.��jN(&�X3W,��#U3����}H�W�%�̴̼�}�b�D]�_���׼'�$t+tBSG��ۉ��y�����8{��u���ʠ;�>�@y鉯H�r���k�_k��� ������Ï�p�N	KB� .�䟄��V9�)�ga��L��� �MGb���%>��-��}m��:�[�E�K�ĈGK\���܉�H�m����ڬ�A�R�˰�ꑩ����y^����"����Ebv#�^"N���H��\�
�!	���]6�W�H��T��ń�.�����S�����&b��
�����B��u��2���T�ӧ/�q�ÇD�;����A!|��4���v�b��S!T��\m$���G"kh�Å���ϵ��a�6��z��Vc��U��j��!M/���ܥ����/B7�oWX�׿�J5X�O2U���"y9������'A`׌懼�\���P(�$g!�+�[����;Jǌ�٬&�I`���NĐtS���n2ݑ������5�_8��^.~���8%��5]~�(�>�NUy���%�O�#w�m��4��\��x����$^v��|l��:?զ��u e������Yg7eݧ)U����S��#�Y�T֨��4&a�q#ljT��4��S}O��������s�y�]�~:6��=@���`>�9�J�U0����>�|I<	W� ,[�/��J�.�?�O�YL=��k��_�V���EF$u��Uz%ԾR}��CwC��y�8b	�`��]e-\�G�x&Qs��&��t9���WZ��"2�m�s���}+ÍX~�%�nfM.��d����E���?��� ],W��D�5�w���lW
���k1�h�ZxPJ�� �J*��_�H#�ǰ�ж4	a�&�^�k���	���������3�L=iI������ψ�r�0P�����-�Jޟ��^��n
�2����zw��^���/���	A˝CdQ	i�'C�,�����WK�E�De/�u���n�JX~S��y��n�K��_W0�|�\�{�%IH>�m˿����2��y��ln%M[���JO��x��|a����)2����/��X�έ�d�qݝ矪Qj�\��3�d���a�����گ�}C-�f�j�����z�,���)��I=���\O�'����?X��L��X+y �����i�l��^�4��	 ��+�~s5Ք�T�p¼������b9�[r��ߗ�s�s4��hCnΨ�	�'D]���Ŭ�"��퐌��el�&�F�����-����T�����aH�n>#u�"�B^�ND�{���"��(F���V���>��3��.���.�?���\��2��kF��D>y�b��=���!�t\5j�Jx��~*��\S��wJ�O��`��xG 7/7�F+��P�����_��h'B����'I×�G��K��8���}4e%,����C9,	# ��&a�9r �s4Ot��E>YfR�i���#Xv}��H��Ef������c�ح�K���"܎9��G���z-@@���p��@�4�ʴ#���Y�C�|M�����H�ޮ��e���;�J�i|vZ�8��p�g$Z�#n�e�ķF�l�Tu�x|d�<�5)��	�#Ã�����Yl����o�Դa��Q,�P�d�q���@2۞9 O�+��O(S�����0�WYF�iO�p0��"{�L��Z`�B����q�B}�H�]6�TN�e.<�$�'��F�ѽs�lf�}�}h�{,d*;W\�VUuÖ����x���r��UZ�"5%Bק�P�}c�w��h~�Ѥ�Qv�6퉆F�^C(�IO�W��̥D�k���F��v�t�U6�#�(��p�ޓ�so�:MB�R��
��;�)�:v.q�ĉ=��ڠ5�b�����X�~��y�J#$LJ�c<q������7�Tw$���V���t�e�מa�=S>���t\h����I�/�Q��?���v�Y&H�RR�w�@TÅ�1S�\'�b~|5�y����g&����b�@4��Y����g�m�d�̾*:�ɮ��x�HZ�|�Em��Nc%���H��W����Wep����S<��7�2�k�$��3���5DqH�D�qqp�����;BA�D3�����-#ï���7�1�kBS)7ɇT����h ���y�]�I*`AT������$�Ё�l�M���7�o�ʁpE[��c�����ϑ�p���Fϭ��{/p[S�%~C�ߴX��P�/(}�y\!ot�8��%��d�b��
�=�h[�_/�Jv�/Oř��W�D�0�΍���A�"�Cl��4����]��u<��ў=k�.nIn� �8���H�r��lϲ���Q��T��d�(bv�,^2��� n� � e�JLgy�+G�^˙f�����m�/h?��)i�ߔc����G���$IqH�<PI�b�H�+�G8���z\�a�O�Nau-c��ﴔ&F�SlN�l;ߤ�@4���|���-�EI��3U������!�ܯ_�h�+y��>��>%V���p=����)̮�e<nl!�����Y*2(�F��	؁^�ڃ}��>+��,�C����Ԡ��hk�n[��/B����5��2o�@O�ګ��1�����u� B�X'��>�,�-�h��Q���P���'�ڊ���=�