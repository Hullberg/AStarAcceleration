��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�Lw��K��i�J��9�P������5�3K���p��	� �!&Ȉ:i��2�����~d~ji-�4	i�OB��Ќ��4RG�	In��%������Ե��!e�ԕш]G�<��w���S|Cwd�L�<s�\
�^�W-z�L�1-X��C%uM�O9�F�H��d����K�B`-��U���A/����u��+�r��%�$'l�~����嬑�X/H����Q�%��˨m�a�] HƴE;��a"���ߦ��C1�F�2Ȉi����7>�^,�s��"�(t�m��ҿ�=<�Z`��Q+<X�A]�D�.-
P5`ax�>��{((�%��p7r�5RWB�!P=#[[����~���=>��U�[�����^�^e���{t�h��;�AzSh�c�ð���_k+��JKI}��Z1lMf�V�i\G]+	��i ��N�Y�"�M5�#�9����u����呰������%�;��{Й�]r���#�7��RJ��c��%��2_�=o��ѯQ��L6���pQ������_X���~�*�H�f$�^^W�YU�@d��4�)��|"��2�C{����r���:�>[�q7y�D<_�-6	�T��`L�g��o#��A���?�S�]������H�5�!~�cB�>O�?�?����a�� �Ş���H�9_���7��g��,��g����׈�'>���m�G���װF�x��b ���p��$�3}������z�An�f�p`	���Uķ6��q��:T�;�~������7�*�9R���E�1j��E�NDWG��2p����N0�����vx��We�N�;v��Z���wô.����Όvխ>[ԩ�P��i��J��.� x��,���+��f�
3����s:�f���׵�����?�����+=��Eg�Ǫ��}s�\QeU|<��*��g���Ӕ���Ȋ!��;��4����9�1S�����a�\��Em�9���\@Və#�m(ϯu��8Vu
1�.\r�e�.	ꦆU"��aIr����5� AVUy"Ct�8E徦K_3���_�����C"�� }��v�����K���ޔ�����i������yK�,�c���j���S��0:ʠ��).B�!a�6�-#�>���I?U|<,������+SI�R1%�q=]��}lq�;Z����q:
���b�$냍X̯P`����(�hW�;����	���tN:���T�D�p�Z�
Z@l|�	v^�/s�EB�Z��dZ82Y��0�У6�0f��r�ӬS����nРR� W���[eC�'�N�T�FuL�F���윟a����5ɢ��
!��}�,���P�hlӃ������S���/��i��?t����N���Y��X� /0�L�p�?a)��E4GDMG8&@-Y��ٙ�,E��8�೐iLo8:=LN�����CL��������t���7b���[�#�m��{�J�`��[DQ�(Ͷ�^�¤T�	�q����zvӁ���Q�{P�-��?#L�/0L����k�d]�{��Ä���X�Q�D���Eٿ1�T��Kh==��m�0��=!9-BA3�@�
�7����!��N�]�R�l��d<��zp�1nbh��"k�H��ۅ)���,"8� C�t�r�C�ZƲ�:�d���.FGۂ��{���1YR�e?N��RJ�d�@��9_��`@�+�@�5�ݢ���KSh���ب�bm/C]�j�R�]ϩ{�GR��x#����D?`"��VɎ t��
�'��1��C[>)����6�Qs&�-J��m0�d0�����˫1wL���A!�5J�z��BިÃ������+�B_��C[���ɩh}+��|2���io�Q�����4��;�тъ��$��B�@�z>�g����7�0�W-�1�|�����Ԋ��������9h�9(����8���(T�a�X`�D�%Y:����Z܆��:ɉm��Z4c�E��vN[t&�֕�h�Q[��ʞw���G�^/利q���q�&���X`;u��=�*0r�a����i��כ�2/���e���'`�����ϲ,`�#�+Eb�ۭ���a-��Cm��O0~������J��)� �(��W[�9�&n���9M�Z���۬|��:#���Vr�*c"Pd�D�u'bFj�>�롺ܷ�&r��_f[w2���Umu�����n��
���	=�����*���c�	ַ���a,��&�����申��1c� �Qj��.�ǟ��[��}h�Y+�r]`���^J��П���Y���s��Y߼�E�1I�J���^�{��IL�/�A��X�c��E���@z~)��ba�EP�>d�0^��0{t�C��h�.T�]ta!�R�%`<�H{#�y�M�@����˕��b5�,l�ȫO����u��)Mm}\1�V��|59�>��-G8�L ��t�x���ތ*�lu��VN�'v�'*bj,`$��	���k��`=Wq�%J@���ǥ��Ox�Q]�X�1Ä$�N>��	�Œ�|I��01��Ѝ�B8�W���w��qT���l2�j1���ɕ�F������wj-Z:��\��X��<��s��Vq���v&��V���YT��|pA� ��{F���R��Y���i*���Y�?�I. ņ8N��Yب�p�Z�o&%T�7��+�oخ�EL����!	�?q����A6`�>�BUA�ל���L<�t���GD�#�ڷC�+۰ն�����UOΚ�