��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���q�����W�E�9 Vοօ�̷�S�;(B�����",�U�s����6���i	t̂9։l7�ڶ\g1?bnL@F���	��;r}�ȓ�d��ٟ�p��p�	�W�E+� ���xp� ����� ���.���%�Cf�Ѽ�#�x�9����T)mLx9�����SCyS<�(6�̍;m��؍�{��<g��((.Z�W�9���+����OJ�:2�	��'�ˌ���{@(��4|�e�$}�~��e�k%���` rE���vm}ӝ;����:1Z$�`Ă�׸k�Ő�J�s��I��+z�#֍[w̢"�\ato_��ӵ��b��W6/Ξ��FG�ϟ=%=��{}�~F�I��|oQK(߼4V{�k��K��'�H�(6L�qk@,d�|�zt�v6�tի9!�@��*��C:���7��kS�[I, [�=�7Xg#d���&|��Hu���Fv��/�.:��?�%n)�ٮxJ��YT�kT�m�OAԾ6�׈��/	���<i��c��� m������$"��^V�>>���A�0�a�HSc-ŕZa�2�~ �D�P��>�Jr�铸�|uXF�(��=A�3�Ucϕh��Y�$!��i7t�4���Qe�����Mr��Ǡ�Z���r4f�P<L�31,��z֦�'��ǟ�U編B���SfW�c�C٢��V�L/�c�conw���3#_�H�{���د��� )���S�U�����E��c��B>ط��n��b�� #��V�ƒ�)ɖ~-�rq�[��,��vQ�$�!bFmM#��Us8��A�4��Ed=f�y��K={:{IϠk+�e[-�p�\ކ%Ǝ�o������?�ї����S�0��	�l�>	nAr��4*�z��EѶ�@�=�`�aX'ڥs{d�5��d�л/�̃Q��8Hˏ��ZP@�Anx$/����9M֦X��U9��������.F����FJ�u��ڳ�I(q�w��!�h�0�Q��J�
K�~���p ���X�(c�d��iJl�y�:�CzpSO��,
�M�u�)J��$�����歐�&�fO@u�}@�h���8����r1�ܨ&���>C~�)b��`f7;��h�L��^"	K6s��bz�a�m"b��-�ϥ�I�(\�nz(˧�/
����0��xm�1~�(�EGN�B����,�42�ĄҰL%�sU�*�����O�V���c�z�z���Oh�b�Hh� mWl�Fn��j"�Ccq	 �M���%nTrR:wM�0r�� %Yv�,&ƭE�1��m�px �C|n��ҹ"� ����F�h��e�g����o�f�Q"׬2cE6��^.|5o�*��Q����]�w��%���<a5�wNGT�U���p�G@5t�����Q�DC����k�04p��'���˃:��X?9$�՜]�hܻi�C�uu�Ι��%�&<���-:�$7a?��Hs���F=�7�|�}95&'�8@�L��8�����k� ��;��@(w�"T|����w\g������/���}�����]�0�5�"JI���h��)�_�2)>V��<Eov�KI{��/���"���6<"G�8����w	e��y���I��_#�V�w�ƞ��i^mf0�Ih
b����:�u���� �y���̊���x<2������VS7N���8d��E��%I3�_%i��Y>*%��K)��X��.���W�A8�ӏi�� ��}�M��"0��C��Cm0�E��V$� ��(�~GL���gAҳ7",��>p�|!���ÿ�`1x&j���>&U>Gp��I!8��u����)�m��gU�=1k��}M\���l��r�U�����&��)TIJ�a���-�1_e�wQ R�u~�N`V�¯iY���"f�S��tq�6�l�}A�-�O�*�~�3a����<��\"c�9��@$�L]�o�l5gw,ӹIL�T��V	����S�b�vB�����E��Abw�������l�^�ZO0�����4� ���7��JG"��9��Ɂ�5�*r� j� ��=����e^_&ˍ�}�M~뼉{T�7�k
�\��>H�.(��10.Lx$�!v��Ώ��0���C_B�4-��ʐ��d�{̍ۿ�in%��x2�#��uJa�k�@"��Sd��[a�kN"�%��������=�b��ϊ����m]��Dot�{"�����>�bj���czs��˚�dKyd�"ýmn9Ϸ�>5��!Ǉ�H%,s�+����Sx�Q��*^89=IΛ�L�Z�5q��$s�z�����ڃo��f֡X-�]����A ��C�Ŀ�8I�����5�p�A��$z9��xm`��<0.�ek�H���̲l\��3C<�N�� ��vɭ��UN��~q�P�A��K��Z-�������#2Xx0b%��I������m�uw��1�ٸ�����Z�����G�k�kv=+V n�?L�	0B����j������ĵP�ܝ8E@�h�*���N�S�ewFX.^�Z�M��:��uw�kk���E}��1�$�At�
��FKf#�q�Ԭ����ݷ��/��2��	��W�]�Z�>L��աf2#r�*Tko�x8�@s#3��0��l���E�ó���w���DK�4�2�5��R��t���"%�Lk̔ܞ:&]�k`�uq2gT3�5ܬ -�
("<x�*�/����ĈP�l�#i��k�u��)o���Hc�]����$rR��/|��ĜR��]�Ղ�6;Rx=rt��� ��n|�<p�Z%P��u�۟�F�qlO`�����DjB�J�xNuL���-�R�˹IM[��eT�W��:�B�k#C�'xNN��6�	�.y8���B$G�,��쑓��F���#��PG������xU�����,e6Fr�?> @Ŧ�r�j�$��G���r�<3�iA����V��G�{D{��~c+����M�yM�n+�٭e>��;��-L2���b(~�ů
���ݘ���4�dr4�T�c��d��r��H���_��