��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸�a�MSa�ĳ1X
�|I\�{pc(���o8��?V�;mN����^2f�����z@���/'
"��$��m����D�jM��'(�}��'\;���gz�F
g��lz��l��H���4�q�
I�}���u��QV��]��� 6	\w/OI"D�j��i���;�O�-j�'�#�c��PC���7�߮�H�go�����o��s�;�x0��J_���ٌ�<���wthG�%�Tg5����mG���߀?m�_��3��x���Tr>%)����ޖ4�.�|��qv�|���P��<��v�;�T� � ��kG�XYPעq�_�<kgl�����������!$�RY���q���r�R=������
�hi�ڼ��V-7���]��U�S5%Ej݀�{RM3п�L��i~����Y6TV��3K8.+�[HJ�e>����'+���Rk?�w�0�;v�9�`D�#R�b'E[eH�>b�M�Q���Rp�p�:O����Gd:|�^2���.9ƪ�V�,چ��*4�����u�A��ӯ�ON̵F�K�Gk[����V������9�`�jjl��W>-�\�P�J���@��Ǡ�|�ś���DmՌ1�~b��,Ø��dƪ��7�����6l�XM�3ϹlBP׌�KׯQ�v�E�?�N��+k���qUR�o�2�����ө�M�>��� "Q%�ﴓu:��Ǣ�W��w��g=�˾ K4����LTT&0~?b0��R	�߳��|��䧜qA�*}EGr�SܤUmo��b�G�ǯT��ci�&��I�-yt%.P=���c�>��x	&[�Z�N����n�m*���ʵ�|�G/�T V�=�S6�ePޅ�]jJ��Ec���l�S;w�AF�T�(��kb?W�c;�nS>��c{��	������w|c?��J��DB7�<�����7��>�����^#)��L��v�&-���מ�-��{A�
�M�<<�A��W�ֳ��(�?���_p��i�� ۻ(|v�f�92�|]�o��%ǽ���Xl�r_H�}^���\��5�x�s���|�P'�wW�D�7�p�� ���������0�櫵�ز��\_���;���	���"��&z�8����J��p�P]Ș��W\�swˆpzB�*v�l.D��٤Q�F��?�u,��S�,/��m��"���IњcwŎ9�`���R�0�N�RK7�������+{zl���)��X�^���J� U"���_ab%��PV��f�*G�h�4$��n��2}P��Oa����YV"u�/�
z�*畝���ť���g�4wZ�o�`��X�%�����ͩ��^�MϠjrZ���y-�Z9�������k!/��'a@��x�%aO��� �Oa�Lϻ�#�:�U����^������+��dȹ^4�ދ.�}Xǚ��g�h�݃���Ǹ�]E�����w��^�.��s��[1�Tn/�$wn�n~5m�Y���K�z���)�H6��&MC *6�Т�$�*6*�����,���^��j��/`�z����ʗ���c}{�ֆ�&Дa��2�	%�8V��9N���owMރˀ�vI���ۋjQ~
�(^8۱`�����1q��f��Okg#gGx�ʪ��&H��������JT�
Xo-��^�#�q��ģ,���3��U�xS12/�:ǎ��7�Bbw�gׯ�(,�1��XMv=�@�u��#��͏�z�M�&1�g5�]��Q�G���J��{�5k�8d��f�o�lH�LL�B�����S���Cˢ�<�f���.ÙP-u��=i6T4�H�����'w�QN5��	t������&GL�Q���c7��>̕���3U��ag�S|:A]>��U�#�-��c�w�z�br/������\[eaю$�@-�fU�P�i�}�{�b���j��9�*��|Q=c�����k[�<3z���[��� 0�T�R�?��F���ɪd'8�Ѣ��_�)�}%����z~D-M� fa�vE�*e���	�
Lή5p	|<4�*�a�j�w�w�چ̖���_���J��dKD�����!�ކq��(�K{Ń��}ص�5S0V�c�-�6q9�s�V���w�1]P�׋R�d��8z�,X�8$Iv.17����U肩<�$�t5�Iv�ǒ\�e�Y~�+�F��g��B�gF�%0��)ߌ�b������P<�Ot��uK��>w�e$=JE��|��I
\���s��쒂I���٪B.\o�M\�D1�mW'��硵G���(��B�H�,l"�<��vT�y�2X�N���@��q��W�x�ȱ��௣�w�lM%����U�iQ}]��jj�'���
�������m����B�689	d�D2oyK9_W��@	�Yj^B�υ����h/YJ�![�����B���������	�Bx�h&��h!w�w���Ҩ���t��cu�M��� ��lw$���=��h����ҼvF>'��5b���xp �H���Ԟ1������Bt�����ph�t��m�vR�˓�CH�#]d�U�9	)�@G,��2��{��Z�m����z�}8���#2{S$��&ȶ<��"�G[pN���r���qx�P�5\����n
0�΃К���xm�^>ṹ}C���C�.���A9KX/��Ǩ��Yd�yB�B�� �p��h�$��Y�Yg����4����Ѯ� %@�k`��.��v���>}�l��ض��Jփ�G�a�l0e����a�9���zUe���Ye����%�b��Ko����	D���@Rϐ��a6l���׌گ��:��>=�+ߠ̯0r�8{��i&,�jeG�$�N�(������p%{ٹ�A�D_��X��zhW� 
��jSwu ��2SJ���a��_�d�N��{�ogGi��t��i8 ��6ݤ��0�6�_l����y���ڏO����������1��YL3lL�7FtU"ñ��	�oh�=m�5����7~ٻ�S˘��gH?�J��tF�Ra��M$��#H$|zͽ��r'q�VK>����L�%�|R��J��ư`'K�0�IO-�0�8��ք� �a������n,7�Y���z�ɲ�I'�C��34������$]I)]
K!��?�47�WO�
Au*�HJ�f�=G������`)�_��v��� Dl���e=S��)\��`۵�&az���z��˙�B#�ov��Up�O��d���d��ײ��x� Y�C�A��e���Z$L��*W��e�O&�7���������SrP�zׂ�U&:-i�T��/x�(íGrg��[�]��mb�|�ݣ�0A��4z���)��E/��|6N����{S�:�!�T�OKBx�)�!���,�$��X�//��$���J�-qI[8ry~�M �1a�.\�+Į�.�[чĊ���@z �n 9u6�R���E<�(#^w�,h�9�~��	��@��^J�'���!��M#�����<��X�(�T���=8h�
�І/��������?��C�$M��>���Xu�jԮ�	>&AX�k�K�n�F�_
ADz��=lMmZ�K��D ����c䨱�:�7 Y�[��|�53Ae��������5u@��/�Mب`�!ӳ�ڴ�ج㼵B�E.��F��@<g�k�