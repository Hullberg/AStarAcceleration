��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���q�����W�E�9 Vοօ�̷�S�;(B�����",�U�s����6���i	t̂9։l\ֿ���Yܼ�^}�N͠y�e��{M�;�L���z=���5!������8�[,T�F��X	����%>��ʦ�a��{fF1�b��Q��_��x�ϥ�@�BB߲�z�aฌ�!!>�P=�͇��m�n�������i8��< �� *�\g�OUE
)ݵ�!�i�
����L�	<�Mi����/��(�Ga��$W{��d,�yt��v(� u��#������Z�UpܨN!�|�vC:�+��'k;�l�S�t��g���5� ��a��;� ��0[;���M{��ȉ��T�]l��4�[:��}nfZ�vP��5~��k�� R�5
�~���F;&M��4�ߵ/�
R���V�[�����>ڸ�Xw�T�d���RE*X�r���;1F�_YiC�̽�~[��(_1��ZI����l貜k���D���F��B�x���|�t���8'Kr��a�G��q��v�\.�>'W�1Z��6�V�����Q�A�7��7,գ7@ˉ�p���z���f�,H<+�|�I�/�6�z����!�e����1��ҝ��t��Yuo��1@9|&����G�I��$��>R{����~h Q�:���ٌ�F� ��:|!w�����O�4��b��s���r�EfB�_pB)(�s��eb�)��Yîd��$��/_8*篗I��D�V3>�	��r�N�Ҝ����&ƍ�й>�!������ǝD��`�^ZU��q����Ә�)l�8��<2:�[�����9꿴9:f��\[�|\���1m(nE�rl��M�� �[j��	�>Mӓ:���saLtb^����d�����K��y�Ǯ�i4�7�n �WHm+��!ڀ�3``l���.P�ɿA,)�ah��ŨV}��pᇢ��x�w!Lkz�y�
��3��5��%q�f�3�Ƒj��ὯC�~�Y`��M؏ ��������њ����*�������K" _Y."��A���N?�$y��|�Σ�^jq��s]r��Nd��/���ߠ�Rٷ��/�AH��mgf���6Sl;w��B���9z��p���r@[#�Ȝ#�>�r�9~YW��D�u��r���˔����s�u$��HL��;*m��٬@N�. �7V��t�	Y��1M��۪�d��Å/�����o���((�=�� a]=v$�]���(ުO&[^}���`��)\�b޷ڒ8a�+f��\�85�q4�������T�12C�ݥ��gB�oջʕ5Y*JP}��9�1j��pNf���H�9z�I$�B����y	֭����X�ZkN��0A_������ S�'ہ�.�Q5X=,d®B!����P�F�����3��:�J����F��X���{������?;�9���ɀܛ��j�����-Mt����������kS#a�h��d���� ����J6�~@[l���4�/��2�O���*-��9DAFKI���-䩏5s���K�߅�(��o@OC�VAe��ؙ�'J���+c������b �=F�ⷔ>
N=�p���6����D���z���Y�S�,J�z0��Da
E|y���b�م���XΧ%b4��&�����g�x9�G��Xi'kpt�A���jr��y��G�9�^��N�ޤ��R�����@��+Խ�`z������K���*�ICa��aR�)-��bR�JA��*��MC��.t�y�/�0k���\�|G�����\�O���u'�X*�UNn@��}������f6Btۨ[f*���@ko�rq�_�<=�$��D��wv+QNꐢ�`�E*I�W�^��y��i�_M��g�s��.Y�k*�3Y�遱���}}O����}��)OMfW ����l�P؃c���r���CE��<Sf19����^�BW\�[�eɱt�x��m�e�R����.�P;� Jr��> ��~��J��ϫ�գzc)����}zQq#�g�Ru�K��ý�D�`�癘>�{�,	,a
��ƕ�T���!1��A�
��;�~�������x�(��b8�qpw�B��J�K��)����8���x�;e�&�ÿe�3I*�+�Ô쒺}��R�/�"����y�l��(7B�Z�}5�꾪
���)���ᮭgӢ,?|��R�"M��2���u>��_;�~zB[LfU��g�deu�3�R1���Y7��.S�Y�sk���&���l���I��W��������0oc��{���q�X�{\:�4���Pօ=�^D�8	A<��Dx@�ޤ#<	j��w��k0��6+�j$�H�^�����3f&��>8�ɏvf�^C��)x:8��p ��1������8�cF/������K[��Qn����W,W��j{ RV�3&�0��kw�h�~/lZB2&{�ă/���+;W��E��9��L@{�7�߻��ym���b�Vvt�(qڑmO����2D���1�D��&�xyTY cܑ1=U<B��\1
�F\6C ����Uޟ	��7<�� �ä	P�6+�v9HW1��3�����G2U���L�w�%�]�ݡ��"H�im�7�o�i�n���H0��~�NF��.�r����@�P8?a�Ę�gZ�l�Z�d+6��ɲ��5㻯i7�\(��:�g�E�H�a	b�)(L �:R`�NZ�L`�6�r�@��Ϻ�&%�[�(/6�(�::<Z�U}<�%�9��E��J2X����R8e�������",nb"�<�|�#|�̵�I���`eT��:(��}�ow@'��*B�,6�T���]J����[4�o;�<b;��H�Bu����\ۃ�γ뙱^�.�Ԍ�]��qi�P�ܾ I05��қ?]h\uu�)�S�����0�:"NR���؊���](�*�uuq��j2�F��dx�E���۸�`E _T�O�񗻣i���˛�Y��z�_u,�y��h�2%�LH��o����Ϙ���*K\��7�7�,��֍M.��1�:/9�� 硏9��A���e%fH�(e��7)0�����F�9ܨQ��P��i	�s���f���]C�#��N�u���E;]T̝�i����݉� /v��k��i���y�����K{"Ic�&�.�u� ���E��`V~�����k����X����yw�S�Z
;��V��"��B�������Ms�,4[����Q��P��Xg�;�^dk�^�����)�U8wy=�	�3{�=�|�	���"����H�����%��6v�(�>ܴ,v��o��j ��}��l�:q�ڈ���O�S��;;t����O�o �9�Ho��/���K�c;N�އ'Br�rk^K�Ö�����%��t[��0:��g^+�D(L>�
��}��=hb��#MO]���n� L������x{]�r���QMwR�V� ӛ��R�����$�贮����[�ZB��k�C�$`":f����k�駏Q�X�F��ߠ����)��1�b�%�Oͧw���v���zE����G<�;[��ނ�)�zt6S�=%D�� kڨ�)�&"Wu�^�6����P�H�[�ֈ���̂3�
v���B8ٛO^�[?�e�����m�Cs)\һ�Na$#���h{����kr
aWX�峳5 Eg�ŀ?Q?�DE@�6�C:�;�<��8�b6MX��UB��8�Ss�Q�X��9��������r_rhV��݄�4#F�C�y�Im��0}�fvCٜF9F�3�!�Ƴ���E��B�t���mJ�u���,o\:^�[��9�����B�I��+=e|m��?c�x//�lk/�+2L��q�3�ő�%A��OdӾ�S&"��n��&,_�֬��8V;�H��Ŵ�2�bj���6}ilˌ��"�.�T��ti,�v��fn\3�[��֗��֧~���n�md1���R�=Cu�X����ނ��JT7���$� �q�zI��+�uf��`ߒ��?�&b���^>|����]=�;h�f�r܅5eŝ�g��>�msY�ߣ�^��9!0�~_2п�� �T`����G��U�ױO���8=�|�8�H_���%`�K9��G�r����Uw(��3c~��R�/�4J�f�B�h2?T�lJ!O�"`+�5�38�2T����H�|׷.�W]��s�9��>�\G�6����e�>���vx�a�B<��Җ�#:�&v�i,a!��\���+Co��F�:�� �E���%�M���ߞZ]��qq����Ww���x���RB�����+�a/�qA-�I�=��1&�|�bq<���L����Z=	�N��)���`�ƙ"uў�����C|q�uu+㒊��m�S� ����^�(�ԅ�у�k�$tIœ|#�