��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸�Σ�HڂͨgT�W�1�.�gW(�CpzQx�E�.�@�6��"o�0_d�hk� 2~!��|Go�E�,�+��ۏ0I�*G�Fnk�#(N�0���w���e�ԃ���D�:�����:��f�p�%9�M1��,^Hg�4zI*w�5��?���Nl�êB�Nzz{*���QӱS� ���Γ�1G���~�^a|���35�t�D�$�8�Y����t�~HgL��(��{��y�T��:�+��W�7��������1�-L�F�ى�*lV�r��-�\��H�x��P[TJ:,����h%��FT����E;�����9��=)�	o
���Eҥ���Z��{B��?cs�����C�%ݚQ�Ӻ�?Fլ�<x�����d͘��_+n�~����L	<�+Kf�Wqd/��3?`t���Y`�<ˉWYzN��<�e�I:"��v�h�lvr"�59kU����l�b%�l�O w�:�-E;��ت@�3�������脇��x����}�(^��7�56s�ے-46R��!����P��`����pN�M��� �"	��Ҕ� Z����z{&[�I��Az�W/�8��@�S
�)�J�R踠����ڬ�zA��dH?{tп����A����c�������=�e�k-���5�e���4���#*4kgl��U��~���\�������9��N)�����3��	6
��9���B�3X��	�Q�]+3E�ș�F�͡Ox��ʠӊ�(�^���H�]�3߀,��^�5W��