��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���i�ƣ��uMdĿ����{&]����W1��d��씒�f�4��f�����¬��g���sK��G�(�'����
��!����[X�~͸���l&ܡf��I�c�w
�Y>���^}����8]�L��;Q���qm,e9��Աuű���z�B׷��!� �7��[T�-�N�v}vk��� �ȕ���2��"H����� ��9�"EB|~�>}5/�ԭ��Z
$��غOGy����{"Z%��m���R�ȍ�#�H�`tq�ѓ�Nc�=���?�`�F��
�3`�"D��~�E��%��o}5p(/f��y�@�B���E��8�}��(3��JG3r=��&K��⋽�IA�����v+�����JGc2)\���;5���T��*�(���̚�[ޗԓƝY0ǍaT�b��t?
_�׏nT���kbT^h=:҉�mP60���ޞH9�]HH��6Ӎ��d*"�i#�&akM��`�i�����>����;̡�֋���W~(��0��/ۿ2(�H&���P�^����Y$�����R�$4�K�3�Ɩ���	���}w��̏ ��)+��A����h������Ȇ)	��R*#lhl3Qz]����.�Ͷ��F��8�Z2�5n:9����J��̉�0Q4���5��ݗ�1c��[Nk,���3���M������TtG�s���U�^.tX蓮��?i��66c�J��b �UOX���}-�I��5�xV?fZ�gg c����_��U�L�y�p辟OkJ��K
4hWn���ܱ(o4X�u<���a;hF�`��Z�^MOFX{c=�@�%��9$	�K��w̼Q��m�l�\��0ͶCqÎ��E��E���zA]{�b�&���"�uOW6e~�撰���|��L56ʿ��-���Q���S�S�'�D�=cw�� 0t1���A����\�NV�S6m��b�z�H�Nn��XK����/8=���k�W/,�����8�i�'�{�����h�<~�0^��P���l����NP�U�/��PeS�h�Lt%6�E�p��Z7�X|�X�����t�{���'r4�I81Fka���P���z��)��׳�����\  ���H�X�5�Rk`��eg�	��g�e��w��Q�M����ddN*ǋ)w��RE���ڄX�A�v�9�&�$�aL�/���ʒXE�	�<����~
w0ϴ���o���� 0!��8|`������RQ��e�|���lx>�@RK�m+uT���JC�j�|�#L��n
sK�	T ��'p��*.��a��O��{���!���Ė$����@6$s�B��������u�A,?���R�=���igcǔX������ ��xY7��ĀH�5A���2"_cxɸ}fC\yXɸ|}���~�3ǃ��LaB=[�[	�cG�*66����c���JLIf~�v�7ބ��Φ)"�P��I˰���e��(���^[��I�u�2�͂f6$�aӶ�������1I\Gӻ�P@�)*���j�Fܲ�M�g�
7} nP�6��]m"�QE]&c\����E�Qw^_-r ,�M�;���&r|�F+r��]�������y��ЇN*�Ɇ���	����g=�%��1[0�����4?����k�b�j��"��/ ��7��U�8+]OQ�6뗸ݭϰ$$��|~�%W(W��N��u-ށ�ej����Rbsw{&\��Ír�ss������lׂ� �#�ZB�n��/)�7����Vd/��y�7��I��fK��~-9�)%�3����.��Xb$�@񴒛�����G���x�HA�"����qR�\0�l�N>R���J�@l]�l�Rs�88�/V?�|��5����a�x�kn������h������eg�f�҂�e���0��Gvzo�"�;	$��
�pqκ,��S�����g��{����p-��R�{�'�^ 4�r$�
��0{l�\u? ���a&��}��o�;&����J+Z�(����'Ѯ��dp_�&��-h�jP�Xq��9�:-W��C�u����|�{�q<��ayк�y݆#:�ik�rx<B�E2��U��P����h�v�C{3�^��+�m.�v��QZ3�1��B��B�++pZ�ȭ_��qZ�D��!�j�$��Ǩ��w|���`�#\"P-_�b�OĎ 6��,�4���"��O���6q(���d�50g��ǟ+ ���D�0�����ג1@���A}��!M>>mt�i8S��A�稬?���$��kv:&�'�qO���&����u�ef�*M-A�;��3����%wDM�R�� ��QXa,�L���Q�ůN7u����XBf���m<�(S��5�e�����=E@�_��#�߄8���i�(w ���Z�s��?eX�L�c���C���Z7�Vz{��QG���[�4��:���5w#Pٻ�\���;Ƣ�Q�F�QKX���[Sе��zL���PK/�H� �g�%"=����H���慕AܾO�+I5^o*Y��'`]��ϓ@�W��;q�C>&>8�ޗ,Rm�y���1�T�Z���+��9���g$O�!�u����v����f�dX���T	1T�#�Ns��#E޹���%��tU�h�[������d�t@9�g���>��W�LY׎3�+��2reJ:�I�1|}%/(cW25��C�i��#e���9�����-1�і���Y��|�l�f�b-c�7�0����;[�V;����i���~z����/��qZ��h��(�X{�z�_wX��Ҕv'	�%`<u�[���������-�S΀WB1Ջ��N-5,��L����I�l��K
��Ǉ��rF���u�"ݓ��dێ3��F��b'B0
��l��>pj���QA��Qϸ���Ez�)�U�uC[y��$���[V,uX���iF�
�(.�d�������<��j*��a��R#��b���*%v��7��h�b�T?�"�XQ��Н|���ll�h�ޕ��#�&���Ĩ'������b}��aN�2�,[_t�&ӆJ����(��A�p�#?;���Wg���:r�m�w�҂\θ �7�I>s��l� ���{��^����#+��E������J<4}�[�>��.���S�y�`$�����
�\4ZT\�y��򋨣��ɿ fk�,� �b��K��֯&��#�	�􁦤98@р"1��"
[����ن��%���B�[�Ed�lͻ�95�1�r0�� r��O9�(&K,S
�b�(�H�
U�Ftc07fV�2Ŭ�=�8K� ��qu���Z[rh����8�0��J�J��_W�ʖ�?H ���^nc��n��&�p8��촬�P��3�l�*�j(��G��(JI	�������c0'kH����g������uM�рI�䥃k�q���nr��L[~\i>K�L��xd���4E�5�y�#�q��kϤ�[͑�MQ\&�+ݹ.�ON=8���~܄.�ЬQ��f6� !��e�ݎ��A	�}Ԗ�4A�rk[�ca�S����&�<��ZI���1c� � wE	�ē��5X��
�}�K�x���.��~ ��NX3&a��}����S���-~��R��0��Y�Kv�vY�K��#4*�/��qh������N�䍻��i��ݗe�h+)�Qh�I�W��{���Qku� ��粹`��nr�B��Jb�K��yZ	�$T|>Ds쨝�-�G]�qNEҸ�|���{��3w�m9���c	�\�,�%��X�����>ejdV�������M��7��g�9�t�C)09X�ĭ�0qbN�ޱ;0�[���}�e7���3_�	��֦�|�"ߨܲ�OTBewP��g��X6�����!zb�Ӈ��N�	��1#�P�>O�"�w�~C8��Y`��U��G�X!<y������k��17��+��D���U�*w�r���r3u+��/�ɏ��V� d����\��p�'�!NT_�
�ۅm&'�Y�7"���նWk�?B��<Ï�q�#��B�F�8VA�׹~��r�&���qy�X3�V� �VM��*�+|r��tbI�sa\Yf����t�aP�S�S�L��T�CT� *�6Y�oΑ��9���L�{�e*�N�~?��?	��Uf���y	".�|���X�����(ѡ͡x}F۫+�!�C�SJ��EX��iA��O��<~&E���.�E����9[��1U��a~�T�tɝ4!?Av4Ӈ�E�Ĩ==�e��2*O������`���\DV���(�>�s��:�^{�Ӹl�p"��M(2Ro����RO/��\B�P[����m�����E}�x/�noTƅ������x$�٫DL)�����A�����w¾���  �5l�*�?�'���� o���ﴄ�%gc�{Zw�.��p�{js���V�ۏ��#�ӆ�#��y����B=z|��T)���o-����3���O;噼���Q��?�_EGE�@Αs=2��0��.���<���-�2GK�,#>�޴�t?��m��z���o��=0��c'��[��b��hw�%�r�F�V���2(#��)��7jziu6�z�DZ�~bz�ס�����e2�J(
�;֚�����l���*r<�܆I�{;��dqPR#�#�S��z�%�*=L���c/h���"��X��U?r�\kL�����{Pv��BZ���՘\{s�e�ת���7�h��X�V>1n�α/�E��B#�cC]�\�Mm�OƗ[]@��CE�eu��b�&����0>�"E<r�L���j��{D���p�����9� 9J|en��7$FM�Ɔ�;������x^��ȋ�T;G����4�l���au�xuշ�#����&-J��a����'��wp������1�Ý{���	M/0BG���?3p]vq��K���f*��9���7���%=]��9�S>(�0RM�j�n���W&���Sd'�{�@4�YT���	i�'��qL�ӕba�vp�~���.�=�4x�G�J�����%9Fv��? h���t����!7��|P* W�ڣ̓1��7�i�T�]���@�X�D��G���gAuʊ�	�o ΃�Կ�^%{0���M?$�jZI�ɉ��fVCK���Zභt�ק���=���]ƠJzI�(g�����
�z�	"��Ö���
1�7��5AI��|�HC��v�f�,��8GtfE��x�EV�L��@3���&S؄���vܩ`��H��wS�s=��3������ Q<�{�.���ƽ�5��u5?�[��W�M���\Ħlyg��фR�Q���]�-d�GV��k�\%�H�E�|Tل��X9���gl�ҕT)�O:�+��Uhs��Zy��`N��6y���]��i�,տh �%䈦ŝ�y��Ca�epʰ(&�с���*�Y+�����K��(��ji<�����\��;���y$�� d�Ȭ����2�<��R�U<�22��ȍ�Vv�ٟ-?ETm^׵0>
#Al��!vg6����q�v�Б�X��CI���̬R7!!`<�{���I�ZJ�
:z��+�s�}�m���~�ަ���Q�B���~:qLr��g���KA�g�R�(�s+B�[޶���A�>�9��<nO��ک����L%ME�xh�m�4��6�;Jr\'��!�[.�-_�������9o�^>�(�v���Aj&J��@[^�V:�}T�x��ӆ[��MyeH�6><w�o����NbJT����7�]�mE�Ÿ�֗�l��E��(��λ�>��D�h`�w��x��մ�%���y�
KO(�\w�O�d�P�B�%@��#�pҞ��ϱ!�hg�i�F��L^OÔ�&s���@����@�<��mW*TE-e�3�p��'�3!�f�Ec���j�}r�� _D���8m�];K�"R�ּ
U|)�GC�̆y|�{�����2uMj��IUxw"_�^`ɀB�ʵ�S��8/�r��+r��e:���j��]$\G��ӡ��p"�A�A|A�+e2I���r|��#%bE�f���F� ���K��M�M��[s��o����Lq[�v$#������q9'i��I���o�G��[�N�p2��1o��l'�?�GF?-a|�yr���OL���s&	�~ˀ��4�������Ϟ�]��F"NCd�/�]�TpCܥ�_\�=j]5"�N
>k�Y��!~���3��j8g��20����fLl=CgA� �x�N�?�VO�dVA`��!�Q w�\@$`ZU�8س#f5�1�sh��LC��`��[.vv�%��x�K׏5}�!CBa�1�Vc�l�H
�����*0]K\��ϝ�H��v)I>j\6�PxO��L磒e�`B�ٽ\�2=g���M�n�hS���\;�<���G��TQ����ZY�K���xKi�)|ۻsFoNO&��He���Iue��� *�E����9b9�r��h�T�K�h�G��������`P��µ|Q*�y�����u�����`i'�:5�
�AJ�S3˔��{ڦ'˱l�x����� ��$�|&���Ӌ}n���_h}.6su��b��i�z�$�BX7,��83 ����@jq�)����Y�c�k�#��E���kf]庖&�(�
B��*д�(Ӈ�U<Ϋ�fH׳|�]���]�ͧ��h��p�j�����0�*����ƭ�8�i}_/�3�L��k��o>:e�M��cq|���i>�,#��T��;Q�����N(o{04`	�h��?��;�;�]�����R�~ډ-�U��<�D ?"���3�<�2�J!I��Y"l�ӕFM�_�`� f��4B䌃�@֚E�5I�׹[Hjս��"��*^�q䌋:�2�	`հ:�i���OQ!��1:�3nϲ*�p���M�?(������86GV�q��j߽Xzz@�B#��ʸ{�����S*8_q�,3h�[��	mz�'VI9��݀��
a��?��'%]0������?R6=�0P� m��`s����˰ptd�6��E&ט\>��%Z�����+�#�d� ��&��T���Y�Ǯ! F�?��Z��
m�Q�j�8�֚��ʩC������X���=�&�>s�Ǣc3�\�����w	��� ��/�e5���o+	�/H��}W�y׵(/���%{ųS3k�Q��ͨ��7��;�<���-|�>�}}�@Ӯ��ّ����M��7(�����n�͛�4�.q�����SҩV0A�LKv��1���!�t��s��!��5�RN�ڮr�l�.e_�-�7����o�M�.�f�N�\��_��0��*A:��������g�[��I���,*�X��/��綢�x��M�mW�,\ȋLJA��������Q��>Čޚ��BY��0���� C��ݵ���W(x���M �WY\ڧkW��S���C m�2��,g��aw8u���|Ն'��Ź+'�Z��8���C�q4�|��\�FA�N��č�	b�Q3�;��X��Vj4�M��T��j7Ʉ_�_?B8򤺊����L;0��>��ea���԰�������{��C~j�1l2�MC��σ�(�����~��
�&��ܪ�.���x�І����d�޵��Q/��pt"49�?׺NN-ҿ�y��*5���9��Dn��Ё>����Ci��!5�
�P��:Pt�3)��Q7A.�7�R莭���i���B�����	���_R��;��L����P��;�V�
Ϛ�{|���r���qs�R������< 	tҥ
�cϨ�����?'kqt�ᬍ��«�5Sn��:�ͼgy�����F�ǎ�]�`��]�Ij�%���禮p���AkE0dπړ��k�^1S&��A�M�:Q0%rq���f�B�
$W�/\l��9��֜j���b<8Q�cy��������H�Q���Th��A�;�n3X4�vSbSIL#�_T{��?֎0g��!�J72~��J��dJ�X�d�ͪXPu�&�Cgup���<�0���:wms�'S��^K\����ԊM��AT:�x<��q�����:�Q6�j��#<I�x��n÷��oA"�2	C=R��w,���8j�^V�/��Ap4Q��$�D��h���78�\3+�j�S���)f�	��N�Cm�%�O	+
� U,'	�0R(Vy�4	?D^z������̯X��[��6��̞�e�6�@�Ê�%}�;��I!�(�ҋӱa����%Հ`$'�P�W��'{����^�+ھ��Ħ��Щ�/	%��!����%T�;�cJF�����\��T�^�����M���rq�S���?:��$�N�x)*	�@z��R����� �{�e�wYZj_�xf��T���xf���g��`���i�j��Q"OrTh����)<T`���?f����,%Շ��l�;;�Rr�w��D���	
�ңiJ:���WG��e��hNKK���e�o��|бR&���1�g'�� �цr�v�{Q���f�|m�)��?ƢE�F��t4�b�$#��lp'7���lZ8K��[=�q&�-~��gB�{�7H��i�͆��f+���A�G�ڗ4���?2B��V.���s� �0$,���+|����-긤�]m~(�\a��??N׳�jX~DB!;���&(���'�� l���6�Iԉ�1�s�?��<�_Z�KR;nAuU�r�B&Q�����N�h����&������j'6M�zNz�^��ʕ2����T�%3��|�'M6�r��vz8���<�i�氡6O�x��!?�:G�Q���:[wb���C��=Нun���W�z/{t@
@���4u���9A�@��V�k�p<��8����سu�`N}	�]i���v�])g%c�b���g<�Jۊ��ۻO���v��I
ߍ>��}X�趼�N�*�%"(R|D)繂A����X4?���:r<�r�
�0��?ƍ�(��8�%��8.6}�Y�AM�/�q@A(#���v�*Ȇ���5<��l���f��8�L4�#jİ�s�?�Ds(��}b��i�]{�	���9ţ��7�?�����B^F�N|�Y_F�x�c��G������'��Sk5o*r��g	�Y�A�1#d����DM���I�P��fgĝ촣���Z���S?ȟ����p�����F.����*�9��+P��J�y�6XV��Z�!~���Z/���Z*�pK�0��t㥼@���gx_�2�+U{�gp���y�c�8̘03�m�H解�coao�g�e����n�������.Ԁ�E�KX�nj��E_��13����6EZB�U�;�M� #��i	�}ͩ�oP��5�TzK
�	=���5m����ݡ���Pq?�qϔ��^ɕ���&�L�#�H���P�$)(���Xqm�Պ��q��I��^�;y��<Ѫ2,_�Ҏ_�ϸq�Fc�6W����x�t��5&`Z�ฝ������x�S�/e�e�"��g҅��![�֗���0(v+p���F��G�ۦ����!�`u����at��'5
INE����㌃%l�b/��c�����)� F�;^9"9����Vq>T�����=�WA��2g�AW!F-�:�2�#^�y���R0/���H�?o�X{�vɠ���b8��ٸT%�kr)q�Ft���Sj����F�>�qS=��d��h	ԆKԶ.d�s��S���N�kg=p۞/E����vdс��brh�;�n��`]bKc�o`@Τ�K�S�H�蹝?�x0;����KV��AY�Ԥu�Eȥ}�@����y�?`5�9lл��-5z��Si��g����	������r]�4�]V�?d`�g_��ȗ����nƛ'>_�h*,bъ)�*�H�`�>CR�r�tpप�1ز�{�<+�Gޒ����&1�	���U��卥�'��8Y���כu�'9�B:Ð�÷	I��������o��;��B[�`U6ג?�;�"�ol�3 �R���f)�r*Yֳ9����ذ���Xi��ۙ
mwm�-�.��B��Q�Z��C�Y��JߌE�`!��A��O��O����1^�,&�`�
S��U��H�B>�6�s)
��?���x�帝jh~��r��O��x�1ci�p.Y�D�V>�W�����wd����?�����!��g��oY����Gp�)Ӯæ������}b�u��AI}��	��8z��k�x��-)V�U�aٜ랜�$C �J��7�3�������.}�M�l,�>�������Wd  a%BΡ6֔OQ���P)k�.��~l y*����g��x΍��ێY�/|��zf�v�~ֽt/�ukc�v"�n���`bq>�T'�b-�����_-��k�������5�J��P�0���)��귽�,��ݒ�q�����A,�Tw�V�^�x��]"��L�'E3lm�R*(��.Y��G�5鬀���3F����S2	�%ĭ�g�g�Tv_�h�.VS'M?p��#���)�hu�?��L��Z�M�^iǭU�=�.���?�tɆ���[N�o=U�����Z" *̺��L�
ɢBl�Po8�IC�_De�B��B���u�a&}.��o�yT[i���d�a���&M
no��Rwh��رO-��ڛw�Y\����w-�	Cr�) x %v?�f����гvDt�Y� nte:�H�J4���C��,'�8}Cx����J���~���R��{d���Sy��+�����Sf��s��g�Z��Q�-�-n��#��	��8E03pJb�|*�̿V�(4۴������W�����˂45	�����[ޞ�J����Z:D	:�B��h�r���E-��?ɋGƯ=���n������b�� 8���ƿ���ڬX+�Αmz�w�F!��75��9qtc	-au�?�.m����۶(�Xp.8�U�
����+��E]�6�O���nw@�t��g�Ģ��-v�֒d�K-���(��4hl�x#i���<�C$�?0��g��J�8y��FL�8H�����XzB�bB��csd�Ӊ��liadLJ��qeh�/'��fZA�oFs*�;�R�g��tJ2mni|o~mX�prMߵ�
��H6se����5���sХkȡӣ�
]w�)��0T��=؟��}RHX>{$GEs2x;c=��'��Pn� �۵=���LLp� �"��A�˵��nv�޻%��aF���X����[��[�̱��:��b��G���!��'S�m�Q�Eﭪ�r��y�j�o�p����Ý�}cA/i0���U	̈́e���Dw�ƹ���/�(�Ե�˗7���.2d�-T���x~�rkRu�;�xKk�:���b�Z-0��3�<��~ش=����)�Dud���H����_`~ï���I����c�ڜ0}�F�M߮��VE��d�C��MwO����~���[L���CDK�ȣƭ��u���Z�+��-`$E�y�L��p���# �ʘ��`�s ��٫C��	��KXr�iV2�U�P��C���raw���W�^��B��I��O�tB	���x\J�[�)�y�j�攻��w���[$��uU~��H�H�� G�<�%�!� ��_;o�Å�FY�c#�C�̏��|��[��'d�N�"�B�6[C�{v*��X�_�?���I���0���胭�FZ�e��E��Tu��[^��\�p+��`|����P��Лb�mR��{^J��~�N���|('N,H�mg�����L�Q�>`������ҧ�ˇy"/� 	��4��������ѣ���c)�2L����I=��5�78W���b�����x����F��
8�� ��(��B���@�;�Ȭ���B��84J�{&{YՖ�q2���t����@>hN����N
��p��ZiW�(�M�{��l��6��]�����2f2*��ݼf� �CM��!D�-�� ���F�Ղ�PR�Py�p��@ ��)�����&��O����,b���)޷@�k'�h��^�po��;�Mv��/�x{ۆ�*D޸�"����c�D�*�g<����������U+e�P���7�%�dp�v֕��D�\�P
K��l
UW�Q�·�R���S@�D�8FV��3!�}�C�c�yl���0�������+��t�b ��
��	�� !��k�%�z���5���<���;ei�a|� 7���*	g*^�A鬚�ĳ� m0�L�h�1h��)%��GEu������ �B�>�_>��".i��w�7^�ҝ��X��I�����|���ݔ��O�q4o4å�B�.d5U�o�7W���ܑ.��j�Q � �*��y��kew�k- ����V+[Uj�*T�J�M<��C9����29��ބ���Bk��K����o/-�����_��.��z���ݬ���?�6��"?�ha��NZ��*�/�{���� "Pf�'|EF��l]#;�B$��ʺ{/)�<+̨7��� T^�	X�U퐠���ݗ��+�ѣ~p4F�ib\����Nʩ�#k�˱S���et0C%�xYo,�ǅ�����9i w�#�؈)`d5�ŏ����ڹ�-&�b��z7p;�ӛB�oM�w���@,C��v���`Rr�z2�"�ݥ,�>#s뚦)�kc;{_�GOP���ؤ�>�ݳ�ܾ��U�P�����"mt�gN��!�����(��a&zi
�Z��9��\�vr��X3��TX$��-`�a��x���$����,^q��@/�qg���ƾ4ސ|�`��5m=�-�f�T���Q�pO7��T���M�EI�,_J|,��U����1ZΛ[~Bw������3Z��Y�H75Ϟ�у
칮�^Ю>}�NA��<�_�:�/�H�(�כ�(_a����I�`���7��}ص.������!��U�9�~�u�EW�(g_Sq��S�x1�'T��<���Q��>����)ٵya�k��.�v��|�z=LIB�@e���Ѩ�{0t��ɂ�O��S%x���"�L��g�n���N�!�_�,hw��Q�Ն���!5{8#Sh7.�}8�b���I�\VX��	�%��Q�KFQ���b�r�m��gJ���*Y9��^b�
�ZA���>w;J��&����;���UB���0eu�Q�A��� UsA,K8��7J�88�[��F��x}�?�[b*E�EX�m���C��;`������C�	ȗ1q����n!
7�M�:<��x�"������tDB����czb��6c�c��Q�����e��^`z�r�}��31�o=���5�:�I����	�-k:w�]�g���T����5�ଂ���eսM{(��ƪ"Փ�M(�|YC<+ 1��Ʌ
�oO���������'���Ӂ9=P����a��0�z�hn��-�O�Lf�oVcq`� ���7�4"uM�A��x_�H�P��q��&I��C���i|c]?5j*�n�Kt�WռG�R5H�R97�g�d�cr�.�\��S�GW���c��O��#� VG�~y�����ۛVz�
�'X2s/QfpgC$�	 8.2E���>��S}��_|��4�Wa@Ԙ+h���ٌ�����$ӺQ���r�>s&D��L�EV������h	.��&�![eFWh8O����֑�����z�S�M�����n���GR�1��{m�D���j��У��:�j�L���ݹ�/�(ܠ �F�Id��Ook L�N�}I���Q��=���0Ϊ�QU��̑r��(�l�.>>�n	w/�:.Đ�RP�_�2g�_+
�b�<��Ч�
�Q����`E
z�($����r�o���`UTK�� ���\�#1�"�:u>U5���Q��"����EC
X��4H��j� ������!1T��7��.���q-UЀ"���F�Q/���vm�-X�P�@�V�	eBj6X����׆�����'��_ٷ�� �<11��HZ������{q�,�8:���v���Ӛ�D�\�SRX�X��4e����Zi��s���ɣ�����q<�C�#G:���r�~�4DL� �T����q�PN�!�1j��œW��+�!��>���&�x0C����ȖI��*���E�k�.c��PŁ���I5O���k����ڴ���	X5v'�?���	=v���0i=��(�'=U��H�� ��^�J(�'�#�M~����]ܨ\���܆�����꭫"� U��\�g��9�T��A7����!�D���Kf��>q֥�,�Yl�+(�C��	�+�?�6���]K6��G0�F��p�������Y!۞D��n��#��zqW�.CA-$[�J���M�1˭M ,�vi�*��Xt�OU���w��j�.��?y�U�@��[���L�j�Ccp@�.����ɪgQ^���'0RK-/$yh���;�i4sL9��
"�L�O]��� +�Ѷ�3;�D�ka�|��kŲ�ͻ�uyqlޣ���g"da$�K�x�h�-BLQ�g|BT�䪮 9�X~�2q͝�3D0�f����S�W֐ԯ��[�|�6�SG3���ޘ���r�v`�dq·
q����f&'S���uz���J��f�1� 	b`��>�� ���4�fK�g3N ����$?ux*�ӓ܂� D��r�=]#��3v��g��a�QrB/K"4n|öZ���f�7'~��<���ރ��2r��96��b!x9�_6�M����f�/ ���N/@������]���N-��+�^���rR���E�a
ž�M���Mm �;t�Rw�1~ͣ(dI5�K�L����Wߋ�C$�OhT����M4�DՃ���<Lʀ��e�%�d�<��|�f��9��k����N�6�W##��2��hBX�!�3�c2>�X���)iB�`}���Ժ�5�"���8'�-;��D�a�wn�=��{�-���ڝi8�I������-Dm-�z3N�@�[��3�S|mSܮ��lV��^Z9�!�j~��-��t���,?J�;�O!F�cp,u�k����� ���`�߭U):���r��~�/��/�6L������c�
1�9��h�������&}i�aG�Q^PXpI��&�Z�gum����ʿ)9���(6#Vy��1�����G��뼫� �U���T�0�K���MjO����/}V��SX}��� ��%u!kn��m�$z8�+�O�¸ZU��r����8lD|��b����pU&_%2�ً�J���ƃHK�}ٳj]ᱼ�N=�ek�T�鴡8a_��j�J���#d��ǉD��e<N-�dm~�'A]���Bx���u��ϝ�1�nG�C�yP��&�(�a� ��U�� �+'"q��m<^<o��w3�2���;�{��	�5
�4w��f:h�%���6,oe���,N�-�I�t:/c�0n�o���oب3蚝�v���A裤�8��\���L��鞥N��G)�p�f��*�6�:�rSY�ޭ���� ��˴��Kn��VO���no:��L�V"�X�[�K� �8}���D���lOF�f=�N�[��D�m�l�JC�ELLn��@�7�;#'��_b��s�F	\70ź�e��]V=R3��7A���;E��y];��v���ʫ>.���nRk�#�u�zj���
�t$�q��/V�D�mޤ����e
�؛Z�.ֻ�k*��J�ґޥIU;�$!]i����
[�@W�L������}����ʧ0
�I�?�9��v��wq�v�]8wF����$���D�zF�<��2^b��'�Ä�aҍ���2e���Yr�i�>6���GY����_�����'�v/E���۬�{w�O����RUC{D�
"�|�m��q��Gb	r�M�Z����v��N/���淏��,��@���y������"��i&��|B K�((>�¸��W�c�Se?�I%�̌����JX�لᙕe��Ӱ1��&�9K���u��v�M#J��*}�N�B�9eys�}Qڌ5g�ؿ�F��"�s뀮�;ulx]@rƓ�)@D��]���J2탫�a�y�;���h���7Yҍb�� ��^�a�3F�}	v��Cd g뭇l*�}����M�,��^D#.#6m-�r�9�F"ͼ��}������h���5ASP٬�66��`[N�a�.U�H����V Z��>����&�S��q�����Ӓ�UAQ�����ԸCx���ک�{�!��y�	�_����̔qd%�Dg&��OJ_^�ɼ V(y���xs~�T���r6P��O7g o�@"V���{2���w��2�ѵ�SO��h�����1�d^d#��G����g�d�_ �z�彾A���u�pK<�6���sK�ztHWK*����VF֞cR���V�aA\1���*��~?Ɗ�\���'#����}�ڤizjW� ���a���L�z-�}�H�]�7��UgO�mP�KنZԦ��Ҹ�EuT�~k���Hyn�t���	���2V1/��#k?�p;��
|2'G�Ɗ�&}9�R	<�U'Q<8�.Pv����^�3���5��-��ܹSɰ�g���E�!k-�IJ��&%&�X��������bP����kq����jS��A1̰l1g:TJ�{�7�<\'ZGǾ'D����5���A��B��6eq����. 6��G������DSX?3���Jc.3��?-	�-! �W�:��(�mp��)=���m�^��G�W_��˕��s��(�?'@;l��P�Z�[���{[#�K��H�N�\���R�`�� 8��| u�R��i�*˖{j�#�Z �zU�S��o���F�K}��[��8��h�9��v�ϯ2x6�o���!h�|�]L�8����� +&���ˢ)����o�T��Nc#����p}(
J�*X~C)���3��n����xq�*9+��6�w��V/O��W��Yh��o�&[��@���f}��I� <y�p�ʯ�j����,���҃��)�![�/8��of���I��_�ӿ���jlJ4��I ��pO����1�����\�km��ڛGՙ#��G���z�W�:2_�΅Lh6��f�~�6�n
wsH ���&���c*�{��df�o/f��t�fᠻ1 D4��T��4�׾|�_թ��b/jV���]t��vcp%��'�˿Q&&T*�4,{���d���A�W=�Js�b�W�vJ�%F����Ϝ+��+��- ��*8�sR��A>e;]��z��W��R���$=����V.�y�x�"�=o_f�\��g�(�3�	���L��*A1�;|':v0NK �"�Y!��َ�{�C'4�C��^�-lG�<	>Ć����� �|�q[U��C�fL���5&�� �^�O�� �P{t{�>Dd=�q��1������W���X/�cm
e�"�D<=��u�g1#���&�X��U��>�h��Ũ���	������
�{W�h$��f��Mx½��Z��;�R Z%�W�Oy4#�Mx\�Ռ䋲��s���ѐ(�;��Mb�B��ec/;�I�I	r�mf��+��۟��߿hJ9� ��3��lhm�E����k���sPι}C�����v`�����ȥ�8�tH^0q�k@X�\� !��ڭ=]���tq�Ö�Z�5�uNko��Q�z��(;&�l��������?��@���Ҧf K�ָ��=wGԩ�uvZՍ�f�(�H��4�2eS��Pj���Y����҆N+n�cR��+)�=*�ҏ��*�i:���G�ӭ7��9��k�t�O�R��߻��c�m�TFW�dC�rr�X�Ƈ��3�9�S�Ei$���x�ş���27D~w�նw}��Hs;��>z�PܔO[�H~��I��EDcPT�V��~�M�&���:�-���^Uj��5�#�~Cעߢ)�k�_���yb�9�<rO�A��~p1p���<5���宷r��v2"U෉�C'V�@�%��1�r-�:(���"�<�����r�a��r�fN��`߬�6�D�����\����Q+��O�ߊ�]
����#춝d�=`�+��
Y!�+�aHr=�H#E7��\�;��-�4h%#�Fp�s+S6u�Y�?9�6�_�܉N�z��uA�m *�54q���/L$!b'n�{��)��(%3_�Q�.� %NM,��9���$O�}d�:\~F:ޠ̎�¯Ƽ�Z���W�%�ӇF<�7>n��^��:�{�G��;�R��rp�ʉ�̥�zQ���/�v!>�3�X~3�V���ϖvƌ7�f�3�E��"�������S��%�k��M0�{(� ��V�\p���,�3���������tK�2��~P`��vzD�Eɺ�;��c�:�K�6ʌ5p�l1Lx}$��!�j�ˉ(�k�ysZ���yQm�)^3دl�Mq����s���s�<�4��
ʸ
dz[I�+���'���i�E$�7����H<�M��A#_�k��z.��(���{����m
��i(��Wi�����r���eV�:��s�Ʌv�L2�ץ��ư`�J&�ۻ͜�ޔ��a��aW7�i���PW��[�88:	��Q&#lѳ�b�hg���I���^u4P6�͌k}�i��F;ݷ�#�<�ت�[�'��p�{��96Os �%�Hz�6�S����:�l�IBC�ӏ�zd3H��.��aq��rCBi�Y���`���]�x@��S#y}	j���z�N�(\��^#2�2.�kđE~�}�/�T�p�_��tvL,I=�a��l�
��U�.��=Io: _���A��ō�����1��b�R#v��u���)*LQ9�;6����/,3nr�nhr�+�\ ½�6U��1�EC��Ɣ�n��>J�c�����WO߈c~�Y ��Ց�@P�*�-U��F��ڴEy~E�|�N�̵��q�u��(���)R�mv��#�D���L�q4p1��6�{�v|�h	����k�x�.ؗ'J #��z8���xmn�I�荕�:���H���@�|YQy���j��(���6�9Ҙs��R�n�e�J{�J�4KV�G��?P�D�G���ryP��蕌���<$�G����<�/�g+*&G�q�Q �M=Ũ=��ˠ0v��7��z>��Ji���i�p1/�&r���B�$���:뜣�45ZN���a^D���k��So_��U�qa�2xs��Q]?R2Lgjx-��z�Uqyb���<R�d,HD��F�*���:+��z�o�ʅ�	�z3&�t�V~!P�B�9u�x�x�Z�5yb�����}��$L�D2�2�D��B���>+���bn�6&=�Pi�iw��6�i:+�u:�{�d�d �RȽ��$�vz4�d^��ln�t����2����q�P��'�,fCv�b)ۉ�D��S���}��(����l;�N�]�+�~��T�2T���&�)%�}
�Xe"%����|�ղ(B�Ij����c�Va�P����>�'-!S|Ā�5F����d�yb9����~�`��\��@>
��D9WE�����q̈́VQ�#���F�[k����CV��A��Y%TN�p���p^�1���̙�yIY���(,,�;����p��YJ�W��o��l�z�8L�}N���:�o�_K�>B��[��%�CSn��N�^:Y?*#F��[�� (a\���T?���U�Q��!Vk����$�ئkd,*�s�$��^�8F�5h��{�y�؁�Tm�=�{S���W���a� C�%c���p6�I��T���@���!���yfp�`뫃��5�����C���6��Q�R���(� [�X